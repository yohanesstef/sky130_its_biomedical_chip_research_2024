magic
tech sky130A
magscale 1 2
timestamp 1729792052
<< error_p >>
rect -29 -127 29 -121
rect -29 -161 -17 -127
rect -29 -167 29 -161
<< nmos >>
rect -18 -89 18 151
<< ndiff >>
rect -76 139 -18 151
rect -76 -77 -64 139
rect -30 -77 -18 139
rect -76 -89 -18 -77
rect 18 139 76 151
rect 18 -77 30 139
rect 64 -77 76 139
rect 18 -89 76 -77
<< ndiffc >>
rect -64 -77 -30 139
rect 30 -77 64 139
<< poly >>
rect -18 151 18 177
rect -18 -111 18 -89
rect -33 -127 33 -111
rect -33 -161 -17 -127
rect 17 -161 33 -127
rect -33 -177 33 -161
<< polycont >>
rect -17 -161 17 -127
<< locali >>
rect -64 139 -30 155
rect -64 -93 -30 -77
rect 30 139 64 155
rect 30 -93 64 -77
rect -33 -161 -17 -127
rect 17 -161 33 -127
<< viali >>
rect -64 -77 -30 139
rect 30 -77 64 139
rect -17 -161 17 -127
<< metal1 >>
rect -70 139 -24 151
rect -70 -77 -64 139
rect -30 -77 -24 139
rect -70 -89 -24 -77
rect 24 139 70 151
rect 24 -77 30 139
rect 64 -77 70 139
rect 24 -89 70 -77
rect -29 -127 29 -121
rect -29 -161 -17 -127
rect 17 -161 29 -127
rect -29 -167 29 -161
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.2 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
