magic
tech sky130A
magscale 1 2
timestamp 1730019635
<< error_p >>
rect 76 207 134 213
rect 76 173 88 207
rect 76 167 134 173
rect -134 -173 -76 -167
rect -134 -207 -122 -173
rect -134 -213 -76 -207
<< nwell >>
rect -8 188 218 226
rect -218 -188 218 188
rect -218 -226 8 -188
<< pmos >>
rect -120 -126 -90 126
rect 90 -126 120 126
<< pdiff >>
rect -182 114 -120 126
rect -182 -114 -170 114
rect -136 -114 -120 114
rect -182 -126 -120 -114
rect -90 114 -28 126
rect -90 -114 -74 114
rect -40 -114 -28 114
rect -90 -126 -28 -114
rect 28 114 90 126
rect 28 -114 40 114
rect 74 -114 90 114
rect 28 -126 90 -114
rect 120 114 182 126
rect 120 -114 136 114
rect 170 -114 182 114
rect 120 -126 182 -114
<< pdiffc >>
rect -170 -114 -136 114
rect -74 -114 -40 114
rect 40 -114 74 114
rect 136 -114 170 114
<< poly >>
rect 72 207 138 223
rect 72 173 88 207
rect 122 173 138 207
rect 72 157 138 173
rect -120 126 -90 152
rect 90 126 120 157
rect -120 -157 -90 -126
rect 90 -152 120 -126
rect -138 -173 -72 -157
rect -138 -207 -122 -173
rect -88 -207 -72 -173
rect -138 -223 -72 -207
<< polycont >>
rect 88 173 122 207
rect -122 -207 -88 -173
<< locali >>
rect 72 173 88 207
rect 122 173 138 207
rect -170 114 -136 130
rect -170 -130 -136 -114
rect -74 114 -40 130
rect -74 -130 -40 -114
rect 40 114 74 130
rect 40 -130 74 -114
rect 136 114 170 130
rect 136 -130 170 -114
rect -138 -207 -122 -173
rect -88 -207 -72 -173
<< viali >>
rect 88 173 122 207
rect -170 -114 -136 114
rect -74 -114 -40 114
rect 40 -114 74 114
rect 136 -114 170 114
rect -122 -207 -88 -173
<< metal1 >>
rect 76 207 134 213
rect 76 173 88 207
rect 122 173 134 207
rect 76 167 134 173
rect -176 114 -130 126
rect -176 -114 -170 114
rect -136 -114 -130 114
rect -176 -126 -130 -114
rect -80 114 -34 126
rect -80 -114 -74 114
rect -40 -114 -34 114
rect -80 -126 -34 -114
rect 34 114 80 126
rect 34 -114 40 114
rect 74 -114 80 114
rect 34 -126 80 -114
rect 130 114 176 126
rect 130 -114 136 114
rect 170 -114 176 114
rect 130 -126 176 -114
rect -134 -173 -76 -167
rect -134 -207 -122 -173
rect -88 -207 -76 -173
rect -134 -213 -76 -207
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
