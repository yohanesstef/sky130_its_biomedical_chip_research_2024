magic
tech sky130A
magscale 1 2
timestamp 1730527170
<< nmos >>
rect -15 -281 15 219
<< ndiff >>
rect -73 207 -15 219
rect -73 -269 -61 207
rect -27 -269 -15 207
rect -73 -281 -15 -269
rect 15 207 73 219
rect 15 -269 27 207
rect 61 -269 73 207
rect 15 -281 73 -269
<< ndiffc >>
rect -61 -269 -27 207
rect 27 -269 61 207
<< poly >>
rect -33 291 33 307
rect -33 257 -17 291
rect 17 257 33 291
rect -33 241 33 257
rect -15 219 15 241
rect -15 -307 15 -281
<< polycont >>
rect -17 257 17 291
<< locali >>
rect -33 257 -17 291
rect 17 257 33 291
rect -61 207 -27 223
rect -61 -285 -27 -269
rect 27 207 61 223
rect 27 -285 61 -269
<< viali >>
rect -61 -269 -27 207
rect 27 -269 61 207
<< metal1 >>
rect -67 207 -21 219
rect -67 -269 -61 207
rect -27 -269 -21 207
rect -67 -281 -21 -269
rect 21 207 67 219
rect 21 -269 27 207
rect 61 -269 67 207
rect 21 -281 67 -269
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 1 diffcov 100 polycov 80 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
