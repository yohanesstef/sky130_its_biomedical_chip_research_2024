magic
tech sky130A
magscale 1 2
timestamp 1730269282
<< psubdiff >>
rect -80 237 -20 271
rect 382 237 442 271
rect -80 211 -46 237
rect -80 -400 -46 -374
rect 408 211 442 237
rect 408 -400 442 -374
rect -80 -434 -20 -400
rect 382 -434 442 -400
<< psubdiffcont >>
rect -20 237 382 271
rect -80 -374 -46 211
rect 408 -374 442 211
rect -20 -434 382 -400
<< locali >>
rect -80 237 -20 271
rect 382 237 442 271
rect -80 211 -46 237
rect -80 -400 -46 -374
rect 408 211 442 237
rect 408 -400 442 -374
rect -80 -434 -20 -400
rect 382 -434 442 -400
<< viali >>
rect -80 46 -46 106
rect 155 -434 207 -400
<< metal1 >>
rect 48 146 114 206
rect -86 106 -40 118
rect -86 46 -80 106
rect -46 46 11 106
rect 63 46 73 106
rect -86 34 -40 46
rect 102 34 260 118
rect 14 -44 310 2
rect 14 -270 60 -44
rect 338 -119 384 118
rect 248 -165 384 -119
rect 102 -209 260 -197
rect 102 -269 155 -209
rect 207 -269 260 -209
rect 302 -223 348 -197
rect 102 -281 260 -269
rect 48 -369 114 -309
rect 155 -394 207 -281
rect 143 -400 219 -394
rect 143 -434 155 -400
rect 207 -434 219 -400
rect 143 -440 219 -434
<< via1 >>
rect 11 46 63 106
rect 155 -269 207 -209
<< metal2 >>
rect 11 106 63 116
rect 11 -55 63 46
rect 11 -108 207 -55
rect 155 -209 207 -108
rect 155 -279 207 -269
use sky130_fd_pr__nfet_01v8_7XSGLL  sky130_fd_pr__nfet_01v8_7XSGLL_0
timestamp 1730023415
transform 1 0 81 0 -1 -270
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_7XSGLL  sky130_fd_pr__nfet_01v8_7XSGLL_1
timestamp 1730023415
transform 1 0 81 0 1 107
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_7XSGLL  sky130_fd_pr__nfet_01v8_7XSGLL_2
timestamp 1730023415
transform 1 0 281 0 -1 45
box -73 -99 73 99
use sky130_fd_pr__nfet_01v8_7XSGLL  sky130_fd_pr__nfet_01v8_7XSGLL_3
timestamp 1730023415
transform 1 0 281 0 1 -208
box -73 -99 73 99
<< labels >>
flabel metal1 -20 84 -20 84 0 FreeSans 160 0 0 0 DVSS
port 0 nsew
flabel metal1 356 -56 356 -56 0 FreeSans 160 0 0 0 drain2
port 2 nsew
flabel metal1 326 -204 326 -204 0 FreeSans 160 0 0 0 preOut
port 3 nsew
flabel metal1 80 -366 80 -366 0 FreeSans 160 0 0 0 rst
port 4 nsew
flabel metal1 76 200 76 200 0 FreeSans 160 0 0 0 vin
port 5 nsew
flabel metal1 170 -27 170 -26 0 FreeSans 160 0 0 0 drain1
port 6 nsew
<< end >>
