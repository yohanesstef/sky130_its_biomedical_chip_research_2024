magic
tech sky130A
magscale 1 2
timestamp 1730474680
<< nwell >>
rect -214 -348 214 314
<< pmos >>
rect -120 -286 120 214
<< pdiff >>
rect -178 202 -120 214
rect -178 -274 -166 202
rect -132 -274 -120 202
rect -178 -286 -120 -274
rect 120 202 178 214
rect 120 -274 132 202
rect 166 -274 178 202
rect 120 -286 178 -274
<< pdiffc >>
rect -166 -274 -132 202
rect 132 -274 166 202
<< poly >>
rect -120 295 120 311
rect -120 261 -104 295
rect 104 261 120 295
rect -120 214 120 261
rect -120 -312 120 -286
<< polycont >>
rect -104 261 104 295
<< locali >>
rect -120 261 -104 295
rect 104 261 120 295
rect -166 202 -132 218
rect -166 -290 -132 -274
rect 132 202 166 218
rect 132 -290 166 -274
<< viali >>
rect -104 261 104 295
rect -166 -274 -132 202
rect 132 -274 166 202
<< metal1 >>
rect -116 295 116 301
rect -116 261 -104 295
rect 104 261 116 295
rect -116 255 116 261
rect -172 202 -126 214
rect -172 -274 -166 202
rect -132 -274 -126 202
rect -172 -286 -126 -274
rect 126 202 172 214
rect 126 -274 132 202
rect 166 -274 172 202
rect 126 -286 172 -274
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
