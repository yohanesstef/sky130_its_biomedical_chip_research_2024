VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO freq_psc
  CLASS BLOCK ;
  FOREIGN freq_psc ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.190 BY 110.910 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 98.160 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 98.160 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END clk
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END out
  PIN psc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 106.910 32.570 110.910 ;
    END
  END psc[0]
  PIN psc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END psc[10]
  PIN psc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END psc[11]
  PIN psc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END psc[12]
  PIN psc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END psc[13]
  PIN psc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END psc[14]
  PIN psc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END psc[15]
  PIN psc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 96.190 30.640 100.190 31.240 ;
    END
  END psc[16]
  PIN psc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 37.440 100.190 38.040 ;
    END
  END psc[17]
  PIN psc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 34.040 100.190 34.640 ;
    END
  END psc[18]
  PIN psc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 96.190 44.240 100.190 44.840 ;
    END
  END psc[19]
  PIN psc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END psc[1]
  PIN psc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 40.840 100.190 41.440 ;
    END
  END psc[20]
  PIN psc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 54.440 100.190 55.040 ;
    END
  END psc[21]
  PIN psc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 51.040 100.190 51.640 ;
    END
  END psc[22]
  PIN psc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 47.640 100.190 48.240 ;
    END
  END psc[23]
  PIN psc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 61.240 100.190 61.840 ;
    END
  END psc[24]
  PIN psc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 64.640 100.190 65.240 ;
    END
  END psc[25]
  PIN psc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 71.440 100.190 72.040 ;
    END
  END psc[26]
  PIN psc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 96.190 68.040 100.190 68.640 ;
    END
  END psc[27]
  PIN psc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 64.490 106.910 64.770 110.910 ;
    END
  END psc[28]
  PIN psc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.150 106.910 74.430 110.910 ;
    END
  END psc[29]
  PIN psc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 106.910 29.350 110.910 ;
    END
  END psc[2]
  PIN psc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 67.710 106.910 67.990 110.910 ;
    END
  END psc[30]
  PIN psc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 70.930 106.910 71.210 110.910 ;
    END
  END psc[31]
  PIN psc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END psc[3]
  PIN psc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END psc[4]
  PIN psc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END psc[5]
  PIN psc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END psc[6]
  PIN psc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END psc[7]
  PIN psc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END psc[8]
  PIN psc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END psc[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 94.490 98.005 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 98.005 ;
      LAYER met1 ;
        RECT 4.210 10.640 94.600 103.660 ;
      LAYER met2 ;
        RECT 4.230 106.630 28.790 107.170 ;
        RECT 29.630 106.630 32.010 107.170 ;
        RECT 32.850 106.630 64.210 107.170 ;
        RECT 65.050 106.630 67.430 107.170 ;
        RECT 68.270 106.630 70.650 107.170 ;
        RECT 71.490 106.630 73.870 107.170 ;
        RECT 74.710 106.630 93.290 107.170 ;
        RECT 4.230 4.280 93.290 106.630 ;
        RECT 4.230 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 93.290 4.280 ;
      LAYER met3 ;
        RECT 3.990 92.840 96.190 98.085 ;
        RECT 4.400 91.440 96.190 92.840 ;
        RECT 3.990 89.440 96.190 91.440 ;
        RECT 4.400 88.040 96.190 89.440 ;
        RECT 3.990 79.240 96.190 88.040 ;
        RECT 4.400 77.840 96.190 79.240 ;
        RECT 3.990 75.840 96.190 77.840 ;
        RECT 4.400 74.440 96.190 75.840 ;
        RECT 3.990 72.440 96.190 74.440 ;
        RECT 4.400 71.040 95.790 72.440 ;
        RECT 3.990 69.040 96.190 71.040 ;
        RECT 3.990 67.640 95.790 69.040 ;
        RECT 3.990 65.640 96.190 67.640 ;
        RECT 4.400 64.240 95.790 65.640 ;
        RECT 3.990 62.240 96.190 64.240 ;
        RECT 4.400 60.840 95.790 62.240 ;
        RECT 3.990 58.840 96.190 60.840 ;
        RECT 4.400 57.440 96.190 58.840 ;
        RECT 3.990 55.440 96.190 57.440 ;
        RECT 3.990 54.040 95.790 55.440 ;
        RECT 3.990 52.040 96.190 54.040 ;
        RECT 4.400 50.640 95.790 52.040 ;
        RECT 3.990 48.640 96.190 50.640 ;
        RECT 4.400 47.240 95.790 48.640 ;
        RECT 3.990 45.240 96.190 47.240 ;
        RECT 4.400 43.840 95.790 45.240 ;
        RECT 3.990 41.840 96.190 43.840 ;
        RECT 4.400 40.440 95.790 41.840 ;
        RECT 3.990 38.440 96.190 40.440 ;
        RECT 4.400 37.040 95.790 38.440 ;
        RECT 3.990 35.040 96.190 37.040 ;
        RECT 3.990 33.640 95.790 35.040 ;
        RECT 3.990 31.640 96.190 33.640 ;
        RECT 3.990 30.240 95.790 31.640 ;
        RECT 3.990 10.715 96.190 30.240 ;
  END
END freq_psc
END LIBRARY

