* NGSPICE file created from freq_psc.ext - technology: sky130A

.subckt freq_psc_8_bit VGND VPWR clk out
+psc[0] psc[1] psc[2] psc[3] psc[4] psc[5] psc[6] psc[7] rst
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_062_ psc_cnt\[1\] net2 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__nand2b_1
XFILLER_9_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_114_ clknet_1_1__leaf_clk _002_ _010_ VGND VGND VPWR VPWR psc_cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_061_ net2 psc_cnt\[1\] VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__and2b_1
X_113_ clknet_1_1__leaf_clk _001_ _009_ VGND VGND VPWR VPWR psc_cnt\[1\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput10 net10 VGND VGND VPWR VPWR out sky130_fd_sc_hd__buf_2
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_8_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_060_ net9 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__inv_2
X_112_ clknet_1_1__leaf_clk _000_ _008_ VGND VGND VPWR VPWR psc_cnt\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_12_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_111_ net9 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__inv_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload0 clknet_1_1__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_6_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_110_ net9 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_7_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_099_ _052_ _053_ _043_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__and3b_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_098_ psc_cnt\[5\] _050_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__or2_1
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_3_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_097_ psc_cnt\[5\] psc_cnt\[4\] _048_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_11_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_096_ _050_ _051_ _043_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and3b_1
X_079_ psc_cnt\[4\] _020_ _036_ _037_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__o2111a_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_095_ psc_cnt\[4\] _048_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__or2_1
X_078_ net6 _019_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_094_ psc_cnt\[4\] psc_cnt\[3\] _046_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__and3_1
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ net6 _019_ psc_cnt\[4\] _020_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_093_ _048_ _049_ _043_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_3_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 psc[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_076_ psc_cnt\[4\] _020_ net6 _019_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__o2bb2a_1
X_059_ psc_cnt\[2\] VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 psc[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_092_ psc_cnt\[3\] _046_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__or2_1
XFILLER_1_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_058_ net5 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__inv_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_075_ _032_ _033_ _034_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_0_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 psc[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_091_ psc_cnt\[3\] _046_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and2_1
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_074_ psc_cnt\[6\] net7 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_057_ psc_cnt\[5\] VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_109_ net9 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
Xinput4 psc[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_090_ _046_ _047_ _043_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__and3b_1
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_073_ psc_cnt\[7\] net8 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__nand2b_1
X_056_ net13 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__inv_2
X_108_ net9 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 psc[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_072_ net8 psc_cnt\[7\] VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_10_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_107_ net9 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_071_ net7 psc_cnt\[6\] VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nand2b_1
XFILLER_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 psc[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
X_106_ net9 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_070_ _025_ _026_ _027_ _029_ _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a41o_1
Xinput7 psc[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_105_ net9 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 psc[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_104_ net9 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 net12 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ clknet_1_0__leaf_clk _017_ _016_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
X_103_ _018_ _054_ _043_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__a21boi_1
XTAP_TAPCELL_ROW_4_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 net10 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlygate4sd3_1
X_102_ _043_ _054_ _055_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and3_1
Xhold2 rst VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ psc_cnt\[6\] _052_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__or2_1
Xhold3 psc_cnt\[7\] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_100_ psc_cnt\[6\] _052_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_6_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_089_ _021_ _045_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nand2_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ psc_cnt\[2\] psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__and3_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_087_ _043_ _044_ _045_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_1_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_1_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_069_ _026_ _027_ _028_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_085_ psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__or2_1
X_068_ net3 _021_ _028_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__a21oi_1
X_067_ psc_cnt\[3\] net4 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and2b_1
XFILLER_9_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_084_ psc_cnt\[0\] _043_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_119_ clknet_1_0__leaf_clk _007_ _015_ VGND VGND VPWR VPWR psc_cnt\[7\] sky130_fd_sc_hd__dfrtp_1
X_083_ net11 _043_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_5_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_066_ net4 psc_cnt\[3\] VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_8_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_118_ clknet_1_0__leaf_clk _006_ _014_ VGND VGND VPWR VPWR psc_cnt\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_065_ net3 psc_cnt\[2\] VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nand2b_1
X_082_ _031_ _040_ _042_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a21oi_4
X_117_ clknet_1_0__leaf_clk _005_ _013_ VGND VGND VPWR VPWR psc_cnt\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_081_ _036_ _038_ _039_ _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__a31o_1
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_064_ _023_ _024_ _022_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_5_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_116_ clknet_1_0__leaf_clk _004_ _012_ VGND VGND VPWR VPWR psc_cnt\[4\] sky130_fd_sc_hd__dfrtp_1
X_063_ psc_cnt\[0\] net1 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__nand2b_1
X_080_ _032_ _033_ _034_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__a21boi_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_115_ clknet_1_1__leaf_clk _003_ _011_ VGND VGND VPWR VPWR psc_cnt\[3\] sky130_fd_sc_hd__dfrtp_1
.ends

