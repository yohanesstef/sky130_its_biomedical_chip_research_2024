* NGSPICE file created from freq_psc.ext - technology: sky130A

.subckt freq_psc VGND VPWR clk out psc[0] psc[1] psc[2] psc[3] psc[4] psc[5] psc[6] psc[7] psc[8] psc[9] psc[10] psc[11]
+psc[12] psc[13] psc[14] psc[15] psc[16] psc[17] psc[18] psc[19] psc[20] psc[21] psc[22] psc[23] psc[24] psc[25] psc[26]
+psc[27] psc[28] psc[29] psc[30] psc[31] rst

X_294_ _118_ _120_ _122_ _101_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__a211o_1
X_501_ clknet_2_2__leaf_clk _021_ _061_ VGND VGND VPWR VPWR psc_cnt\[29\] sky130_fd_sc_hd__dfrtp_1
X_432_ psc_cnt\[28\] _230_ _231_ net44 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__o211a_1
X_363_ psc_cnt\[6\] _184_ VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__or2_1
XFILLER_3_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_415_ net35 _218_ _220_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__and3_1
X_346_ psc_cnt\[0\] net35 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and2b_1
XFILLER_12_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_277_ net2 _079_ net32 _080_ _104_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__a221oi_1
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_329_ _066_ net17 _091_ net18 VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__o22a_1
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_33 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ _121_ _103_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__and2b_1
X_500_ clknet_2_2__leaf_clk _020_ _060_ VGND VGND VPWR VPWR psc_cnt\[28\] sky130_fd_sc_hd__dfrtp_1
X_431_ psc_cnt\[28\] _230_ VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__nand2_1
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_362_ _184_ _182_ net38 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and3b_1
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_276_ net3 _078_ net2 _079_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__o22a_1
X_345_ net59 net35 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__xnor2_1
X_414_ _214_ _219_ VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_259_ net12 VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__inv_2
X_328_ _069_ net13 _156_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_292_ _104_ _105_ _107_ _108_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__o22a_1
X_361_ _179_ _183_ VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__and2_1
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_430_ _230_ net37 _228_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__and3b_1
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_275_ psc_cnt\[11\] net3 VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__and2b_1
X_413_ psc_cnt\[22\] psc_cnt\[21\] psc_cnt\[20\] VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__and3_1
X_344_ _123_ _164_ _172_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__a21oi_4
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_327_ psc_cnt\[28\] net21 VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__and2b_1
X_258_ net23 VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__inv_2
XFILLER_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_291_ _103_ _105_ _106_ _119_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__and4_1
XPHY_EDGE_ROW_15_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_360_ psc_cnt\[5\] psc_cnt\[4\] VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__and2_1
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_489_ clknet_2_1__leaf_clk _008_ _049_ VGND VGND VPWR VPWR psc_cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_0_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_274_ _097_ _098_ _099_ _102_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__and4_1
X_412_ psc_cnt\[21\] _216_ psc_cnt\[22\] VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__a21o_1
XFILLER_5_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_343_ _171_ _169_ _166_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__or3_4
XFILLER_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_326_ _094_ net22 net21 _093_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__o22a_1
X_257_ net26 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__inv_2
XFILLER_18_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_309_ _136_ _137_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__nor2_1
XFILLER_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput34 net34 VGND VGND VPWR VPWR out sky130_fd_sc_hd__buf_2
XFILLER_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ psc_cnt\[8\] _082_ _083_ psc_cnt\[7\] _108_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o221a_1
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_488_ clknet_2_1__leaf_clk _007_ _048_ VGND VGND VPWR VPWR psc_cnt\[16\] sky130_fd_sc_hd__dfrtp_1
X_273_ _077_ net4 _096_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__a21oi_1
X_411_ psc_cnt\[21\] _216_ _217_ net35 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__o211a_1
XFILLER_5_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_342_ _162_ _135_ _158_ _170_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__and4b_1
X_325_ _152_ net47 VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__nor2_1
X_256_ net27 VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__inv_2
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_2
X_308_ net19 psc_cnt\[26\] VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__and2b_1
XFILLER_1_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_239_ psc_cnt\[20\] VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_487_ clknet_2_2__leaf_clk _006_ _047_ VGND VGND VPWR VPWR psc_cnt\[15\] sky130_fd_sc_hd__dfrtp_1
X_272_ _097_ _100_ _096_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__a21oi_1
X_410_ psc_cnt\[21\] _216_ VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__nand2_1
X_341_ _132_ _159_ _144_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__o21ba_1
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_324_ _151_ _148_ _150_ _147_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__or4_4
X_255_ net28 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__inv_2
XFILLER_13_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_4
X_238_ net14 VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__inv_2
XFILLER_1_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_307_ net20 psc_cnt\[27\] VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_10_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_486_ clknet_2_2__leaf_clk _005_ _046_ VGND VGND VPWR VPWR psc_cnt\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_271_ _099_ _098_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__nand2b_1
X_340_ _161_ _167_ _168_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__o21ai_1
XFILLER_23_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_469_ net41 VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__inv_2
X_323_ _094_ net22 VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__and2_1
X_254_ net29 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__inv_2
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clknet_2_3__leaf_clk VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__clkinv_2
X_237_ net15 VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__inv_2
X_306_ _067_ psc_cnt\[22\] _131_ _133_ _134_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__a2111o_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_485_ clknet_2_2__leaf_clk _004_ _045_ VGND VGND VPWR VPWR psc_cnt\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_270_ net5 _076_ _077_ net4 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_20_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_468_ net41 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__inv_2
X_399_ psc_cnt\[17\] _208_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__or2_1
XFILLER_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_322_ psc_cnt\[30\] net24 VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__and2b_1
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_253_ net30 VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ net14 psc_cnt\[21\] VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__and2b_1
X_236_ psc_cnt\[24\] VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__inv_2
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_484_ clknet_2_3__leaf_clk _003_ _044_ VGND VGND VPWR VPWR psc_cnt\[12\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_3_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_467_ net41 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__inv_2
X_398_ psc_cnt\[17\] psc_cnt\[16\] _205_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__and3_1
XFILLER_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_321_ psc_cnt\[31\] net25 VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__and2b_1
X_252_ net31 VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 net33 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_2
X_304_ net13 psc_cnt\[20\] VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__and2b_1
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_483_ clknet_2_3__leaf_clk _002_ _043_ VGND VGND VPWR VPWR psc_cnt\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_16_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_466_ net41 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__inv_2
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_397_ _208_ net36 _207_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__and3b_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_251_ psc_cnt\[8\] VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__inv_2
X_320_ _147_ net45 VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__nor2_1
XFILLER_1_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout41 net33 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_4
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_449_ net42 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__inv_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_303_ _067_ psc_cnt\[22\] _131_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__a21o_1
Xhold17 net34 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_19_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_482_ clknet_2_3__leaf_clk _001_ _042_ VGND VGND VPWR VPWR psc_cnt\[10\] sky130_fd_sc_hd__dfrtp_1
X_465_ net41 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__inv_2
X_396_ psc_cnt\[16\] _205_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__and2_1
XFILLER_2_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_250_ psc_cnt\[9\] VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__inv_2
Xfanout42 net33 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_448_ net42 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__inv_2
X_379_ psc_cnt\[11\] _195_ VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__or2_1
XFILLER_24_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_302_ net16 psc_cnt\[23\] VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__and2b_1
XFILLER_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_481_ clknet_2_3__leaf_clk _031_ _041_ VGND VGND VPWR VPWR psc_cnt\[9\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_464_ net39 VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__inv_2
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_395_ psc_cnt\[16\] _205_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__or2_1
X_378_ _195_ _194_ net38 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__and3b_1
X_447_ net42 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_0_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_301_ psc_cnt\[16\] _073_ _127_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__o21a_1
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_480_ clknet_2_3__leaf_clk _030_ _040_ VGND VGND VPWR VPWR psc_cnt\[8\] sky130_fd_sc_hd__dfrtp_1
X_394_ _205_ net37 _206_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and3b_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_463_ net39 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_377_ psc_cnt\[10\] _188_ _192_ VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__and3_1
X_446_ net42 VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__inv_2
XFILLER_13_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_300_ _072_ psc_cnt\[17\] VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__or2_1
X_429_ _205_ _222_ _229_ VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__and3_1
Xinput1 psc[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_393_ _074_ _203_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__nand2_1
X_462_ net39 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_13_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_376_ psc_cnt\[10\] _193_ VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__or2_1
X_445_ net42 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__inv_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_428_ psc_cnt\[24\] psc_cnt\[25\] psc_cnt\[26\] psc_cnt\[27\] VGND VGND VPWR VPWR
+ _229_ sky130_fd_sc_hd__and4_1
X_359_ psc_cnt\[4\] _179_ psc_cnt\[5\] VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__a21o_1
Xinput2 psc[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_392_ psc_cnt\[13\] psc_cnt\[12\] _197_ _204_ VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__and4_2
X_461_ net39 VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout35 _173_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_6
X_375_ _193_ _191_ net38 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and3b_1
X_444_ net41 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_3_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_427_ psc_cnt\[25\] psc_cnt\[26\] _225_ psc_cnt\[27\] VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__a31o_1
X_358_ net36 _180_ _181_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and3_1
Xinput3 psc[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ _115_ _116_ _117_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_22_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_391_ _074_ _075_ VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__nor2_1
X_460_ net39 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__inv_2
XFILLER_4_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout36 _173_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_6
X_374_ _188_ _192_ VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__and2_1
X_443_ net40 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__inv_2
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 psc[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_288_ _083_ psc_cnt\[7\] _084_ psc_cnt\[6\] VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__a22o_1
X_357_ psc_cnt\[4\] _179_ VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__nand2_1
X_426_ _092_ _226_ _227_ net44 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__o211a_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_10_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_409_ _216_ net35 _215_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and3b_1
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_390_ net44 _202_ _203_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__and3_1
Xfanout37 _173_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_6
XFILLER_13_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_373_ _080_ _081_ VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__nor2_1
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_442_ net40 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 psc[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_287_ _084_ psc_cnt\[6\] _085_ psc_cnt\[5\] VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__o22a_1
X_356_ psc_cnt\[4\] _179_ VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__or2_1
X_425_ _092_ _226_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__nand2_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_408_ psc_cnt\[20\] _205_ _213_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__and3_1
XFILLER_24_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_339_ _152_ net46 _155_ _150_ _149_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_25_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput30 psc[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout38 _173_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_6
X_372_ _080_ _190_ VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__nand2_1
X_441_ net40 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_14_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_355_ _179_ net36 _178_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and3b_1
X_286_ _113_ _114_ _109_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__a21o_1
X_424_ psc_cnt\[25\] _225_ _226_ net44 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__o211a_1
Xinput6 psc[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ net6 _075_ net5 _076_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__a22oi_1
X_407_ psc_cnt\[20\] _214_ VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__or2_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_338_ _141_ _143_ _158_ _139_ _138_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_25_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput31 psc[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
XFILLER_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput20 psc[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_371_ net38 _189_ _190_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__and3_1
XFILLER_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_440_ net39 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
Xfanout39 net33 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_4
XFILLER_24_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_23_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_354_ psc_cnt\[3\] psc_cnt\[2\] psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _179_
+ sky130_fd_sc_hd__and4_1
X_285_ psc_cnt\[4\] _086_ _087_ psc_cnt\[3\] VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__o22a_1
X_423_ psc_cnt\[25\] _225_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__nand2_1
Xinput7 psc[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_268_ net7 _074_ net6 _075_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__o22a_1
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_406_ _214_ net35 _212_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__and3b_1
X_337_ _163_ _165_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__and2_1
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput32 psc[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput21 psc[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 psc[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_10_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_370_ psc_cnt\[8\] _188_ VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__nand2_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_499_ clknet_2_2__leaf_clk _019_ _059_ VGND VGND VPWR VPWR psc_cnt\[27\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_284_ _110_ _111_ _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__a21o_1
X_353_ psc_cnt\[2\] psc_cnt\[1\] psc_cnt\[0\] psc_cnt\[3\] VGND VGND VPWR VPWR _178_
+ sky130_fd_sc_hd__a31o_1
X_422_ _225_ net35 _224_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__and3b_1
Xinput8 psc[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_267_ net7 _074_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__and2_1
X_405_ _205_ _213_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__and2_1
X_336_ _127_ _128_ _129_ _125_ _124_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__a32o_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_319_ net24 psc_cnt\[30\] VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__and2b_1
Xinput22 psc[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput33 rst VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_1
Xinput11 psc[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_498_ clknet_2_2__leaf_clk _018_ _058_ VGND VGND VPWR VPWR psc_cnt\[26\] sky130_fd_sc_hd__dfrtp_1
X_421_ psc_cnt\[24\] _205_ _222_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__and3_1
X_352_ net35 _176_ _177_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__and3_1
X_283_ _087_ psc_cnt\[3\] _088_ psc_cnt\[2\] VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__a22o_1
Xinput9 psc[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_266_ net39 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
X_404_ psc_cnt\[19\] psc_cnt\[18\] psc_cnt\[17\] psc_cnt\[16\] VGND VGND VPWR VPWR
+ _213_ sky130_fd_sc_hd__and4_1
X_335_ _128_ _129_ _130_ _163_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__and4b_1
XFILLER_2_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ psc_cnt\[10\] VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__inv_2
X_318_ net25 psc_cnt\[31\] VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__and2b_1
Xinput23 psc[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 psc[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_497_ clknet_2_2__leaf_clk _017_ _057_ VGND VGND VPWR VPWR psc_cnt\[25\] sky130_fd_sc_hd__dfrtp_2
XFILLER_24_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_351_ psc_cnt\[2\] psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__nand3_1
X_282_ _088_ psc_cnt\[2\] _089_ psc_cnt\[1\] VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__o22a_1
X_420_ psc_cnt\[24\] _223_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__or2_1
XFILLER_25_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_403_ _070_ _211_ VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__nand2_1
X_334_ _146_ _154_ _160_ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__and3b_1
X_265_ net43 VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__inv_2
XFILLER_2_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_248_ psc_cnt\[11\] VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__inv_2
Xinput24 psc[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput13 psc[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_317_ _135_ _141_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__or3_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_496_ clknet_2_1__leaf_clk _016_ _056_ VGND VGND VPWR VPWR psc_cnt\[24\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_17_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ psc_cnt\[1\] psc_cnt\[0\] psc_cnt\[2\] VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__a21o_1
X_281_ _089_ psc_cnt\[1\] _090_ psc_cnt\[0\] VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__a211o_1
X_479_ clknet_2_3__leaf_clk _029_ _039_ VGND VGND VPWR VPWR psc_cnt\[7\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_2_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_264_ psc_cnt\[29\] VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__inv_2
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_402_ psc_cnt\[18\] _209_ _211_ net36 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o211a_1
X_333_ _141_ _142_ _143_ _161_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__or4_4
X_247_ psc_cnt\[12\] VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__inv_2
Xinput25 psc[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput14 psc[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_316_ _142_ _143_ _144_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__or3_1
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_495_ clknet_2_0__leaf_clk _015_ _055_ VGND VGND VPWR VPWR psc_cnt\[23\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ _085_ psc_cnt\[5\] psc_cnt\[4\] _086_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__a22o_1
X_478_ clknet_2_3__leaf_clk _028_ _038_ VGND VGND VPWR VPWR psc_cnt\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ psc_cnt\[28\] VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__inv_2
X_332_ _152_ _156_ _153_ _155_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__or4b_4
X_401_ psc_cnt\[18\] _209_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__nand2_1
XFILLER_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_246_ psc_cnt\[13\] VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__inv_2
Xinput15 psc[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_315_ psc_cnt\[23\] net16 VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__and2b_1
Xinput26 psc[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_494_ clknet_2_0__leaf_clk _014_ _054_ VGND VGND VPWR VPWR psc_cnt\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_14_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_477_ clknet_2_1__leaf_clk _027_ _037_ VGND VGND VPWR VPWR psc_cnt\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262_ psc_cnt\[26\] VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__inv_2
X_400_ _209_ _210_ net36 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__and3b_1
X_331_ _155_ _157_ _158_ _159_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_19_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_245_ psc_cnt\[14\] VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__inv_2
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput16 psc[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_314_ psc_cnt\[25\] net18 VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__and2b_1
Xinput27 psc[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_22_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_493_ clknet_2_0__leaf_clk _013_ _053_ VGND VGND VPWR VPWR psc_cnt\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_476_ clknet_2_1__leaf_clk _026_ _036_ VGND VGND VPWR VPWR psc_cnt\[4\] sky130_fd_sc_hd__dfrtp_1
X_330_ _067_ psc_cnt\[22\] _068_ psc_cnt\[21\] VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__o22a_1
X_261_ psc_cnt\[25\] VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__inv_2
X_459_ net39 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_244_ psc_cnt\[15\] VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__inv_2
Xinput28 psc[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
X_313_ psc_cnt\[24\] net17 VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__and2b_1
Xinput17 psc[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone2 _173_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_9_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_492_ clknet_2_0__leaf_clk _012_ _052_ VGND VGND VPWR VPWR psc_cnt\[20\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_14_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_475_ clknet_2_1__leaf_clk _025_ _035_ VGND VGND VPWR VPWR psc_cnt\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_25_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ net1 VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__inv_2
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_389_ psc_cnt\[14\] _201_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__nand2_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_458_ net39 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput29 psc[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
X_243_ net8 VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__inv_2
X_312_ _136_ _137_ _139_ _140_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__or4_1
Xinput18 psc[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_491_ clknet_2_0__leaf_clk _010_ _051_ VGND VGND VPWR VPWR psc_cnt\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_474_ clknet_2_1__leaf_clk _022_ _034_ VGND VGND VPWR VPWR psc_cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_388_ psc_cnt\[14\] _201_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__or2_1
X_457_ net40 VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__inv_2
X_311_ psc_cnt\[26\] net19 VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__and2b_1
Xinput19 psc[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_11_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_242_ net9 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__inv_2
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_490_ clknet_2_0__leaf_clk _009_ _050_ VGND VGND VPWR VPWR psc_cnt\[18\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_5_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_473_ clknet_2_1__leaf_clk _011_ _033_ VGND VGND VPWR VPWR psc_cnt\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_387_ _201_ net37 _200_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and3b_1
XFILLER_15_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_456_ net40 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__inv_2
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_310_ psc_cnt\[27\] net20 VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__and2b_1
X_439_ _095_ _235_ net44 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a21boi_1
X_241_ net10 VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__inv_2
XFILLER_22_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_472_ clknet_2_1__leaf_clk _000_ _032_ VGND VGND VPWR VPWR psc_cnt\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_386_ psc_cnt\[13\] psc_cnt\[12\] _197_ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__and3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_455_ net40 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__inv_2
XFILLER_14_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_240_ psc_cnt\[19\] VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__inv_2
X_438_ net37 _234_ _235_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__and3_1
Xrebuffer1 psc_cnt\[31\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd1_1
X_369_ psc_cnt\[8\] _188_ VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__or2_1
XFILLER_6_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_471_ net39 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__inv_2
XFILLER_25_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_385_ psc_cnt\[13\] _198_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__or2_1
X_454_ net41 VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_437_ psc_cnt\[30\] _233_ VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__nand2_1
X_368_ _188_ _187_ net38 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__and3b_1
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_299_ _072_ psc_cnt\[17\] psc_cnt\[16\] _073_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__a22o_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_470_ net41 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__inv_2
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_453_ net41 VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__inv_2
X_384_ _198_ _199_ net38 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_15_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_436_ psc_cnt\[30\] _233_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__or2_1
Xrebuffer3 _148_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_367_ psc_cnt\[7\] psc_cnt\[6\] _179_ _183_ VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__and4_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_298_ _124_ _125_ _126_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__and3b_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_419_ _223_ net35 _221_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__and3b_1
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_452_ net41 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__inv_2
X_383_ psc_cnt\[12\] _197_ VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_18_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_435_ _233_ net37 _232_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__and3b_1
Xrebuffer4 _153_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd1_1
X_366_ psc_cnt\[6\] _179_ _183_ psc_cnt\[7\] VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__a31o_1
XFILLER_13_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_504_ clknet_2_0__leaf_clk _065_ _064_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfrtp_1
X_297_ _071_ psc_cnt\[18\] VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__or2_1
XFILLER_6_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_349_ net35 _174_ _175_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_418_ _205_ _222_ VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__and2_1
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_382_ psc_cnt\[12\] _197_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_451_ net42 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_24_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ clknet_2_2__leaf_clk _024_ _063_ VGND VGND VPWR VPWR psc_cnt\[31\] sky130_fd_sc_hd__dfrtp_1
X_434_ psc_cnt\[28\] psc_cnt\[29\] _230_ VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__and3_1
X_365_ net38 _185_ _186_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and3_1
XFILLER_13_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_296_ net11 _070_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__nand2_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrebuffer5 _153_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_279_ net32 _080_ _081_ net31 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__nand2_1
X_417_ psc_cnt\[23\] _213_ _219_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_8_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_381_ _197_ net38 _196_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__and3b_1
X_450_ net42 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__inv_2
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_24_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_502_ clknet_2_2__leaf_clk _023_ _062_ VGND VGND VPWR VPWR psc_cnt\[30\] sky130_fd_sc_hd__dfrtp_1
X_433_ _094_ _231_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__nand2_1
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_364_ psc_cnt\[6\] _184_ VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__nand2_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_295_ net11 _070_ _071_ psc_cnt\[18\] VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_12_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_278_ _105_ _106_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__nand2_1
X_347_ psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__or2_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_416_ _205_ _213_ _219_ psc_cnt\[23\] VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_24_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_380_ psc_cnt\[11\] psc_cnt\[10\] _188_ _192_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__and4_1
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
.ends

