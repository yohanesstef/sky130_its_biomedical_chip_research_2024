magic
tech sky130A
magscale 1 2
timestamp 1730306127
<< nwell >>
rect -623 605 -576 659
rect -613 82 -567 160
<< metal1 >>
rect -325 1014 559 1065
rect -532 865 -526 917
rect -474 865 -468 917
rect -325 866 -274 1014
rect -20 793 -10 845
rect 42 793 49 845
rect 508 800 559 1014
rect 521 700 563 734
rect -623 605 -576 659
rect 189 593 199 645
rect 251 593 261 645
rect 453 580 476 598
rect 423 579 476 580
rect -282 526 -230 532
rect -282 468 -230 474
rect -117 516 134 562
rect 415 552 476 579
rect -613 160 -567 381
rect -613 129 -521 160
rect -613 14 -567 129
rect -117 88 -71 516
rect 415 488 461 552
rect -342 42 -71 88
rect -43 441 461 488
rect -43 14 3 441
rect -613 -32 3 14
<< via1 >>
rect -526 865 -474 917
rect -10 793 42 845
rect 199 593 251 645
rect -282 474 -230 526
<< metal2 >>
rect -526 917 -474 923
rect -474 866 42 916
rect -526 859 -474 865
rect -10 845 42 866
rect -10 783 42 793
rect 199 645 251 655
rect 199 526 251 593
rect -288 474 -282 526
rect -230 474 248 526
use ncell_pfd  ncell_pfd_0
timestamp 1730269282
transform 0 -1 195 -1 0 900
box -86 -440 442 271
use pcell_pfd  pcell_pfd_0
timestamp 1730269591
transform -1 0 379 0 1 281
box 482 -341 1076 735
<< labels >>
flabel metal1 -602 644 -602 644 0 FreeSans 160 90 0 0 DVDD
port 0 nsew
flabel metal1 542 720 542 720 0 FreeSans 160 0 0 0 DVSS
port 1 nsew
flabel metal1 438 526 438 526 0 FreeSans 160 90 0 0 preOut
port 2 nsew
flabel metal1 -288 1038 -288 1038 0 FreeSans 160 0 0 0 rst
port 3 nsew
flabel metal2 -118 892 -118 892 0 FreeSans 160 0 0 0 vin
port 4 nsew
<< end >>
