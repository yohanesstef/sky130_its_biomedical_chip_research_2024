magic
tech sky130A
magscale 1 2
timestamp 1729853601
<< error_p >>
rect -29 161 29 167
rect -29 127 -17 161
rect -29 121 29 127
<< pwell >>
rect -214 -299 214 299
<< nmos >>
rect -18 -151 18 89
<< ndiff >>
rect -76 77 -18 89
rect -76 -139 -64 77
rect -30 -139 -18 77
rect -76 -151 -18 -139
rect 18 77 76 89
rect 18 -139 30 77
rect 64 -139 76 77
rect 18 -151 76 -139
<< ndiffc >>
rect -64 -139 -30 77
rect 30 -139 64 77
<< psubdiff >>
rect -178 229 -82 263
rect 82 229 178 263
rect -178 167 -144 229
rect 144 167 178 229
rect -178 -229 -144 -167
rect 144 -229 178 -167
rect -178 -263 -82 -229
rect 82 -263 178 -229
<< psubdiffcont >>
rect -82 229 82 263
rect -178 -167 -144 167
rect 144 -167 178 167
rect -82 -263 82 -229
<< poly >>
rect -33 161 33 177
rect -33 127 -17 161
rect 17 127 33 161
rect -33 111 33 127
rect -18 89 18 111
rect -18 -177 18 -151
<< polycont >>
rect -17 127 17 161
<< locali >>
rect -178 229 -82 263
rect 82 229 178 263
rect -178 167 -144 229
rect 144 167 178 229
rect -33 127 -17 161
rect 17 127 33 161
rect -64 77 -30 93
rect -64 -155 -30 -139
rect 30 77 64 93
rect 30 -155 64 -139
rect -178 -229 -144 -167
rect 144 -229 178 -167
rect -178 -263 -82 -229
rect 82 -263 178 -229
<< viali >>
rect -17 127 17 161
rect -64 -139 -30 77
rect 30 -139 64 77
<< metal1 >>
rect -29 161 29 167
rect -29 127 -17 161
rect 17 127 29 161
rect -29 121 29 127
rect -70 77 -24 89
rect -70 -139 -64 77
rect -30 -139 -24 77
rect -70 -151 -24 -139
rect 24 77 70 89
rect 24 -139 30 77
rect 64 -139 70 77
rect 24 -151 70 -139
<< properties >>
string FIXED_BBOX -161 -246 161 246
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.2 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
