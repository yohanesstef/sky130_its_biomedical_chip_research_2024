VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO freq_psc
  CLASS BLOCK ;
  FOREIGN freq_psc ;
  ORIGIN 0.000 0.000 ;
  SIZE 51.025 BY 61.745 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 49.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 49.200 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END clk
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 47.025 27.240 51.025 27.840 ;
    END
  END out
  PIN psc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END psc[0]
  PIN psc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END psc[1]
  PIN psc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END psc[2]
  PIN psc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 57.745 16.470 61.745 ;
    END
  END psc[3]
  PIN psc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 57.745 26.130 61.745 ;
    END
  END psc[4]
  PIN psc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 57.745 29.350 61.745 ;
    END
  END psc[5]
  PIN psc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 57.745 32.570 61.745 ;
    END
  END psc[6]
  PIN psc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 47.025 34.040 51.025 34.640 ;
    END
  END psc[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 47.025 17.040 51.025 17.640 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 45.270 49.045 ;
      LAYER li1 ;
        RECT 5.520 10.795 45.080 49.045 ;
      LAYER met1 ;
        RECT 4.210 10.640 45.080 49.200 ;
      LAYER met2 ;
        RECT 4.230 57.465 15.910 57.745 ;
        RECT 16.750 57.465 25.570 57.745 ;
        RECT 26.410 57.465 28.790 57.745 ;
        RECT 29.630 57.465 32.010 57.745 ;
        RECT 32.850 57.465 43.610 57.745 ;
        RECT 4.230 10.695 43.610 57.465 ;
      LAYER met3 ;
        RECT 3.990 45.240 47.025 49.125 ;
        RECT 4.400 43.840 47.025 45.240 ;
        RECT 3.990 41.840 47.025 43.840 ;
        RECT 4.400 40.440 47.025 41.840 ;
        RECT 3.990 38.440 47.025 40.440 ;
        RECT 4.400 37.040 47.025 38.440 ;
        RECT 3.990 35.040 47.025 37.040 ;
        RECT 3.990 33.640 46.625 35.040 ;
        RECT 3.990 28.240 47.025 33.640 ;
        RECT 4.400 26.840 46.625 28.240 ;
        RECT 3.990 18.040 47.025 26.840 ;
        RECT 3.990 16.640 46.625 18.040 ;
        RECT 3.990 10.715 47.025 16.640 ;
  END
END freq_psc
END LIBRARY

