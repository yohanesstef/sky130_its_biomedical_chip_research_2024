magic
tech sky130A
magscale 1 2
timestamp 1730019635
<< nwell >>
rect -211 -274 211 274
<< pmos >>
rect -15 -126 15 126
<< pdiff >>
rect -73 114 -15 126
rect -73 -114 -61 114
rect -27 -114 -15 114
rect -73 -126 -15 -114
rect 15 114 73 126
rect 15 -114 27 114
rect 61 -114 73 114
rect 15 -126 73 -114
<< pdiffc >>
rect -61 -114 -27 114
rect 27 -114 61 114
<< nsubdiff >>
rect -175 204 -79 238
rect 79 204 175 238
rect -175 142 -141 204
rect 141 142 175 204
rect -175 -204 -141 -142
rect 141 -204 175 -142
rect -175 -238 -79 -204
rect 79 -238 175 -204
<< nsubdiffcont >>
rect -79 204 79 238
rect -175 -142 -141 142
rect 141 -142 175 142
rect -79 -238 79 -204
<< poly >>
rect -15 126 15 152
rect -15 -152 15 -126
<< locali >>
rect -175 204 -79 238
rect 79 204 175 238
rect -175 142 -141 204
rect 141 142 175 204
rect -61 114 -27 130
rect -61 -130 -27 -114
rect 27 114 61 130
rect 27 -130 61 -114
rect -175 -204 -141 -142
rect 141 -204 175 -142
rect -175 -238 -79 -204
rect 79 -238 175 -204
<< viali >>
rect -61 -114 -27 114
rect 27 -114 61 114
<< metal1 >>
rect -67 114 -21 126
rect -67 -114 -61 114
rect -27 -114 -21 114
rect -67 -126 -21 -114
rect 21 114 67 126
rect 21 -114 27 114
rect 61 -114 67 114
rect 21 -126 67 -114
<< properties >>
string FIXED_BBOX -158 -221 158 221
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
