magic
tech sky130A
magscale 1 2
timestamp 1730021255
<< nwell >>
rect 482 -341 1076 735
<< nsubdiff >>
rect 518 665 578 699
rect 980 665 1040 699
rect 518 639 552 665
rect 518 -271 552 -245
rect 1006 639 1040 665
rect 1006 -271 1040 -245
rect 518 -305 578 -271
rect 980 -305 1040 -271
<< nsubdiffcont >>
rect 578 665 980 699
rect 518 -245 552 639
rect 1006 -245 1040 639
rect 578 -305 980 -271
<< locali >>
rect 518 665 578 699
rect 980 665 1040 699
rect 518 639 552 665
rect 518 -271 552 -245
rect 1006 639 1040 665
rect 1006 -271 1040 -245
rect 518 -305 578 -271
rect 980 -305 1040 -271
<< viali >>
rect 1006 306 1040 534
<< metal1 >>
rect 646 577 712 643
rect 846 577 912 643
rect 612 147 658 306
rect 700 294 858 546
rect 912 534 1046 546
rect 912 306 1006 534
rect 1040 306 1046 534
rect 912 304 1046 306
rect 900 294 1046 304
rect 900 221 946 294
rect 756 175 946 221
rect 756 100 802 175
rect 612 -193 658 -134
rect 700 -152 858 100
rect 900 65 947 100
rect 612 -239 912 -193
use sky130_fd_pr__pfet_01v8_SC63VW  sky130_fd_pr__pfet_01v8_SC63VW_0
timestamp 1730019635
transform -1 0 879 0 1 456
box -109 -224 109 190
use sky130_fd_pr__pfet_01v8_SC63VW  sky130_fd_pr__pfet_01v8_SC63VW_1
timestamp 1730019635
transform -1 0 679 0 1 456
box -109 -224 109 190
use sky130_fd_pr__pfet_01v8_SC63VW  sky130_fd_pr__pfet_01v8_SC63VW_3
timestamp 1730019635
transform 1 0 679 0 1 10
box -109 -224 109 190
use sky130_fd_pr__pfet_01v8_SC63VW  sky130_fd_pr__pfet_01v8_SC63VW_4
timestamp 1730019635
transform 1 0 879 0 -1 -62
box -109 -224 109 190
<< labels >>
flabel metal1 979 438 979 438 0 FreeSans 800 0 0 0 DVDD
port 0 nsew
flabel metal1 854 585 854 585 0 FreeSans 800 0 0 0 VIN
port 1 nsew
flabel metal1 658 584 658 584 0 FreeSans 800 0 0 0 RST
port 2 nsew
flabel metal1 633 235 633 235 0 FreeSans 800 0 0 0 drain1
port 3 nsew
flabel metal1 643 -215 644 -215 0 FreeSans 800 0 0 0 drain2
port 4 nsew
flabel metal1 921 93 921 93 0 FreeSans 800 0 0 0 preout
port 5 nsew
<< end >>
