VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO freq_psc
  CLASS BLOCK ;
  FOREIGN freq_psc ;
  ORIGIN 0.000 0.000 ;
  SIZE 61.860 BY 72.580 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 60.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 60.080 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END clk
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END out
  PIN psc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END psc[0]
  PIN psc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 68.580 45.450 72.580 ;
    END
  END psc[10]
  PIN psc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 68.580 42.230 72.580 ;
    END
  END psc[11]
  PIN psc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 68.580 26.130 72.580 ;
    END
  END psc[12]
  PIN psc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 68.580 29.350 72.580 ;
    END
  END psc[13]
  PIN psc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 68.580 22.910 72.580 ;
    END
  END psc[14]
  PIN psc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 68.580 19.690 72.580 ;
    END
  END psc[15]
  PIN psc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END psc[1]
  PIN psc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END psc[2]
  PIN psc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END psc[3]
  PIN psc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END psc[4]
  PIN psc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END psc[5]
  PIN psc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END psc[6]
  PIN psc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END psc[7]
  PIN psc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 68.580 39.010 72.580 ;
    END
  END psc[8]
  PIN psc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 68.580 35.790 72.580 ;
    END
  END psc[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 57.860 23.840 61.860 24.440 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 56.310 59.925 ;
      LAYER li1 ;
        RECT 5.520 10.795 56.120 59.925 ;
      LAYER met1 ;
        RECT 5.520 10.640 56.120 60.080 ;
      LAYER met2 ;
        RECT 7.000 68.300 19.130 68.580 ;
        RECT 19.970 68.300 22.350 68.580 ;
        RECT 23.190 68.300 25.570 68.580 ;
        RECT 26.410 68.300 28.790 68.580 ;
        RECT 29.630 68.300 35.230 68.580 ;
        RECT 36.070 68.300 38.450 68.580 ;
        RECT 39.290 68.300 41.670 68.580 ;
        RECT 42.510 68.300 44.890 68.580 ;
        RECT 45.730 68.300 54.650 68.580 ;
        RECT 7.000 4.280 54.650 68.300 ;
        RECT 7.000 4.000 15.910 4.280 ;
        RECT 16.750 4.000 19.130 4.280 ;
        RECT 19.970 4.000 22.350 4.280 ;
        RECT 23.190 4.000 25.570 4.280 ;
        RECT 26.410 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 54.650 4.280 ;
      LAYER met3 ;
        RECT 4.000 48.640 57.860 60.005 ;
        RECT 4.400 47.240 57.860 48.640 ;
        RECT 4.000 38.440 57.860 47.240 ;
        RECT 4.400 37.040 57.860 38.440 ;
        RECT 4.000 24.840 57.860 37.040 ;
        RECT 4.000 23.440 57.460 24.840 ;
        RECT 4.000 10.715 57.860 23.440 ;
  END
END freq_psc
END LIBRARY

