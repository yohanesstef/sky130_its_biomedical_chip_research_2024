magic
tech sky130A
magscale 1 2
timestamp 1730520524
<< nmos >>
rect -120 -219 120 281
<< ndiff >>
rect -178 269 -120 281
rect -178 -207 -166 269
rect -132 -207 -120 269
rect -178 -219 -120 -207
rect 120 269 178 281
rect 120 -207 132 269
rect 166 -207 178 269
rect 120 -219 178 -207
<< ndiffc >>
rect -166 -207 -132 269
rect 132 -207 166 269
<< poly >>
rect -120 281 120 307
rect -120 -257 120 -219
rect -120 -291 -104 -257
rect 104 -291 120 -257
rect -120 -307 120 -291
<< polycont >>
rect -104 -291 104 -257
<< locali >>
rect -166 269 -132 285
rect -166 -223 -132 -207
rect 132 269 166 285
rect 132 -223 166 -207
rect -120 -291 -104 -257
rect 104 -291 120 -257
<< viali >>
rect -166 -207 -132 269
rect 132 -207 166 269
rect -52 -291 52 -257
<< metal1 >>
rect -172 269 -126 281
rect -172 -207 -166 269
rect -132 -207 -126 269
rect -172 -219 -126 -207
rect 126 269 172 281
rect 126 -207 132 269
rect 166 -207 172 269
rect 126 -219 172 -207
rect -64 -257 64 -251
rect -64 -291 -52 -257
rect 52 -291 64 -257
rect -64 -297 64 -291
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
