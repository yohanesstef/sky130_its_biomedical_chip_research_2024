magic
tech sky130A
magscale 1 2
timestamp 1729792052
<< error_p >>
rect -29 561 29 567
rect -29 527 -17 561
rect -29 521 29 527
rect -29 -527 29 -521
rect -29 -561 -17 -527
rect -29 -567 29 -561
<< nwell >>
rect -112 -580 112 580
<< pmos >>
rect -18 -480 18 480
<< pdiff >>
rect -76 468 -18 480
rect -76 -468 -64 468
rect -30 -468 -18 468
rect -76 -480 -18 -468
rect 18 468 76 480
rect 18 -468 30 468
rect 64 -468 76 468
rect 18 -480 76 -468
<< pdiffc >>
rect -64 -468 -30 468
rect 30 -468 64 468
<< poly >>
rect -33 561 33 577
rect -33 527 -17 561
rect 17 527 33 561
rect -33 511 33 527
rect -18 480 18 511
rect -18 -511 18 -480
rect -33 -527 33 -511
rect -33 -561 -17 -527
rect 17 -561 33 -527
rect -33 -577 33 -561
<< polycont >>
rect -17 527 17 561
rect -17 -561 17 -527
<< locali >>
rect -33 527 -17 561
rect 17 527 33 561
rect -64 468 -30 484
rect -64 -484 -30 -468
rect 30 468 64 484
rect 30 -484 64 -468
rect -33 -561 -17 -527
rect 17 -561 33 -527
<< viali >>
rect -17 527 17 561
rect -64 -468 -30 468
rect 30 -468 64 468
rect -17 -561 17 -527
<< metal1 >>
rect -29 561 29 567
rect -29 527 -17 561
rect 17 527 29 561
rect -29 521 29 527
rect -70 468 -24 480
rect -70 -468 -64 468
rect -30 -468 -24 468
rect -70 -480 -24 -468
rect 24 468 70 480
rect 24 -468 30 468
rect 64 -468 70 468
rect 24 -480 70 -468
rect -29 -527 29 -521
rect -29 -561 -17 -527
rect 17 -561 29 -527
rect -29 -567 29 -561
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.8 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
