magic
tech sky130A
timestamp 1729792052
<< error_p >>
rect -16 84 16 87
rect -16 67 -10 84
rect -16 64 16 67
rect -16 -67 16 -64
rect -16 -84 -10 -67
rect -16 -87 16 -84
<< nmos >>
rect -18 -48 18 48
<< ndiff >>
rect -47 42 -18 48
rect -47 -42 -41 42
rect -24 -42 -18 42
rect -47 -48 -18 -42
rect 18 42 47 48
rect 18 -42 24 42
rect 41 -42 47 42
rect 18 -48 47 -42
<< ndiffc >>
rect -41 -42 -24 42
rect 24 -42 41 42
<< poly >>
rect -18 84 18 92
rect -18 67 -10 84
rect 10 67 18 84
rect -18 48 18 67
rect -18 -67 18 -48
rect -18 -84 -10 -67
rect 10 -84 18 -67
rect -18 -92 18 -84
<< polycont >>
rect -10 67 10 84
rect -10 -84 10 -67
<< locali >>
rect -18 67 -10 84
rect 10 67 18 84
rect -41 42 -24 50
rect -41 -50 -24 -42
rect 24 42 41 50
rect 24 -50 41 -42
rect -18 -84 -10 -67
rect 10 -84 18 -67
<< viali >>
rect -10 67 10 84
rect -41 -42 -24 42
rect 24 -42 41 42
rect -10 -84 10 -67
<< metal1 >>
rect -16 84 16 87
rect -16 67 -10 84
rect 10 67 16 84
rect -16 64 16 67
rect -44 42 -21 48
rect -44 -42 -41 42
rect -24 -42 -21 42
rect -44 -48 -21 -42
rect 21 42 44 48
rect 21 -42 24 42
rect 41 -42 44 42
rect 21 -48 44 -42
rect -16 -67 16 -64
rect -16 -84 -10 -67
rect 10 -84 16 -67
rect -16 -87 16 -84
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.96 l 0.36 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
