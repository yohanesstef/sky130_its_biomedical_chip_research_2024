magic
tech sky130A
magscale 1 2
timestamp 1730101678
<< viali >>
rect 16681 19465 16715 19499
rect 5641 19397 5675 19431
rect 7757 19397 7791 19431
rect 5917 19329 5951 19363
rect 6101 19329 6135 19363
rect 6193 19329 6227 19363
rect 7389 19329 7423 19363
rect 11253 19329 11287 19363
rect 13277 19329 13311 19363
rect 14197 19329 14231 19363
rect 14289 19329 14323 19363
rect 15117 19329 15151 19363
rect 15945 19329 15979 19363
rect 16221 19329 16255 19363
rect 16497 19329 16531 19363
rect 16865 19329 16899 19363
rect 6377 19261 6411 19295
rect 6653 19261 6687 19295
rect 13001 19261 13035 19295
rect 14473 19261 14507 19295
rect 15393 19261 15427 19295
rect 15485 19261 15519 19295
rect 16129 19193 16163 19227
rect 11161 19125 11195 19159
rect 14381 19125 14415 19159
rect 16313 19125 16347 19159
rect 16497 18921 16531 18955
rect 16129 18853 16163 18887
rect 6837 18785 6871 18819
rect 9965 18785 9999 18819
rect 11805 18785 11839 18819
rect 16037 18785 16071 18819
rect 4629 18717 4663 18751
rect 4721 18717 4755 18751
rect 5089 18717 5123 18751
rect 13737 18717 13771 18751
rect 14197 18717 14231 18751
rect 14473 18717 14507 18751
rect 14841 18717 14875 18751
rect 15393 18717 15427 18751
rect 16258 18717 16292 18751
rect 16405 18717 16439 18751
rect 16681 18717 16715 18751
rect 5365 18649 5399 18683
rect 10241 18649 10275 18683
rect 12081 18649 12115 18683
rect 13829 18649 13863 18683
rect 15301 18649 15335 18683
rect 4905 18581 4939 18615
rect 11713 18581 11747 18615
rect 13553 18581 13587 18615
rect 15761 18581 15795 18615
rect 6469 18377 6503 18411
rect 10793 18377 10827 18411
rect 12081 18377 12115 18411
rect 14289 18377 14323 18411
rect 14765 18377 14799 18411
rect 4629 18309 4663 18343
rect 11897 18309 11931 18343
rect 12817 18309 12851 18343
rect 13645 18309 13679 18343
rect 14565 18309 14599 18343
rect 4261 18241 4295 18275
rect 4353 18241 4387 18275
rect 6561 18241 6595 18275
rect 9413 18241 9447 18275
rect 10517 18241 10551 18275
rect 10701 18241 10735 18275
rect 10977 18241 11011 18275
rect 12357 18241 12391 18275
rect 12725 18241 12759 18275
rect 13001 18241 13035 18275
rect 13461 18241 13495 18275
rect 13737 18241 13771 18275
rect 14105 18241 14139 18275
rect 15209 18241 15243 18275
rect 15393 18241 15427 18275
rect 15761 18241 15795 18275
rect 1409 18173 1443 18207
rect 1685 18173 1719 18207
rect 11253 18173 11287 18207
rect 16129 18173 16163 18207
rect 10701 18105 10735 18139
rect 11161 18105 11195 18139
rect 11529 18105 11563 18139
rect 13001 18105 13035 18139
rect 14933 18105 14967 18139
rect 16405 18105 16439 18139
rect 4169 18037 4203 18071
rect 6101 18037 6135 18071
rect 9505 18037 9539 18071
rect 11897 18037 11931 18071
rect 12265 18037 12299 18071
rect 13369 18037 13403 18071
rect 14749 18037 14783 18071
rect 2605 17833 2639 17867
rect 5181 17833 5215 17867
rect 5365 17833 5399 17867
rect 6653 17833 6687 17867
rect 11069 17833 11103 17867
rect 11437 17833 11471 17867
rect 4537 17765 4571 17799
rect 14933 17765 14967 17799
rect 15577 17765 15611 17799
rect 2697 17697 2731 17731
rect 10793 17697 10827 17731
rect 2789 17629 2823 17663
rect 2973 17629 3007 17663
rect 3157 17629 3191 17663
rect 4445 17629 4479 17663
rect 4629 17629 4663 17663
rect 4905 17629 4939 17663
rect 6285 17629 6319 17663
rect 11345 17629 11379 17663
rect 11529 17629 11563 17663
rect 14289 17629 14323 17663
rect 14933 17629 14967 17663
rect 15209 17629 15243 17663
rect 15301 17629 15335 17663
rect 15393 17629 15427 17663
rect 15577 17629 15611 17663
rect 4721 17561 4755 17595
rect 5089 17561 5123 17595
rect 5333 17561 5367 17595
rect 5549 17561 5583 17595
rect 10517 17561 10551 17595
rect 11037 17561 11071 17595
rect 11253 17561 11287 17595
rect 2421 17493 2455 17527
rect 2973 17493 3007 17527
rect 6653 17493 6687 17527
rect 6837 17493 6871 17527
rect 9045 17493 9079 17527
rect 10885 17493 10919 17527
rect 14197 17493 14231 17527
rect 15117 17493 15151 17527
rect 2237 17289 2271 17323
rect 4077 17289 4111 17323
rect 5825 17289 5859 17323
rect 6193 17289 6227 17323
rect 10517 17289 10551 17323
rect 10701 17289 10735 17323
rect 1685 17221 1719 17255
rect 1901 17221 1935 17255
rect 2605 17221 2639 17255
rect 2973 17221 3007 17255
rect 7113 17221 7147 17255
rect 8861 17221 8895 17255
rect 10333 17221 10367 17255
rect 2145 17153 2179 17187
rect 2421 17153 2455 17187
rect 2697 17153 2731 17187
rect 2845 17153 2879 17187
rect 3065 17153 3099 17187
rect 3203 17153 3237 17187
rect 3709 17153 3743 17187
rect 4169 17153 4203 17187
rect 4445 17153 4479 17187
rect 5733 17153 5767 17187
rect 6009 17153 6043 17187
rect 6837 17153 6871 17187
rect 8953 17153 8987 17187
rect 9597 17153 9631 17187
rect 10149 17153 10183 17187
rect 10609 17153 10643 17187
rect 10793 17153 10827 17187
rect 12909 17153 12943 17187
rect 13185 17153 13219 17187
rect 13369 17153 13403 17187
rect 14381 17153 14415 17187
rect 14473 17153 14507 17187
rect 14657 17153 14691 17187
rect 14749 17153 14783 17187
rect 14841 17153 14875 17187
rect 15025 17153 15059 17187
rect 15117 17153 15151 17187
rect 15577 17153 15611 17187
rect 15853 17153 15887 17187
rect 16037 17153 16071 17187
rect 16221 17153 16255 17187
rect 3433 17085 3467 17119
rect 3617 17085 3651 17119
rect 4537 17085 4571 17119
rect 8585 17085 8619 17119
rect 12725 17085 12759 17119
rect 15669 17085 15703 17119
rect 16129 17085 16163 17119
rect 2053 17017 2087 17051
rect 4353 17017 4387 17051
rect 12541 17017 12575 17051
rect 13001 17017 13035 17051
rect 14657 17017 14691 17051
rect 15301 17017 15335 17051
rect 15761 17017 15795 17051
rect 1869 16949 1903 16983
rect 3341 16949 3375 16983
rect 4261 16949 4295 16983
rect 9873 16949 9907 16983
rect 12725 16949 12759 16983
rect 12817 16949 12851 16983
rect 15393 16949 15427 16983
rect 2513 16745 2547 16779
rect 3065 16745 3099 16779
rect 5457 16745 5491 16779
rect 5641 16745 5675 16779
rect 10425 16745 10459 16779
rect 13737 16745 13771 16779
rect 14565 16745 14599 16779
rect 5733 16677 5767 16711
rect 12265 16677 12299 16711
rect 12449 16677 12483 16711
rect 2421 16609 2455 16643
rect 11897 16609 11931 16643
rect 12909 16609 12943 16643
rect 13277 16609 13311 16643
rect 14381 16609 14415 16643
rect 1777 16541 1811 16575
rect 1961 16541 1995 16575
rect 2642 16541 2676 16575
rect 3433 16541 3467 16575
rect 4445 16541 4479 16575
rect 4629 16541 4663 16575
rect 4813 16541 4847 16575
rect 4905 16541 4939 16575
rect 5181 16541 5215 16575
rect 5917 16541 5951 16575
rect 6377 16541 6411 16575
rect 12081 16541 12115 16575
rect 13461 16541 13495 16575
rect 13553 16541 13587 16575
rect 13829 16541 13863 16575
rect 14289 16541 14323 16575
rect 14933 16541 14967 16575
rect 15485 16541 15519 16575
rect 15761 16541 15795 16575
rect 16129 16541 16163 16575
rect 2789 16473 2823 16507
rect 3249 16473 3283 16507
rect 5273 16473 5307 16507
rect 5489 16473 5523 16507
rect 6561 16473 6595 16507
rect 10609 16473 10643 16507
rect 12449 16473 12483 16507
rect 1869 16405 1903 16439
rect 2145 16405 2179 16439
rect 4629 16405 4663 16439
rect 5089 16405 5123 16439
rect 6009 16405 6043 16439
rect 6101 16405 6135 16439
rect 6285 16405 6319 16439
rect 6745 16405 6779 16439
rect 10241 16405 10275 16439
rect 10409 16405 10443 16439
rect 13001 16405 13035 16439
rect 13185 16405 13219 16439
rect 16129 16405 16163 16439
rect 8125 16201 8159 16235
rect 12725 16201 12759 16235
rect 14749 16201 14783 16235
rect 15761 16201 15795 16235
rect 2053 16133 2087 16167
rect 4997 16133 5031 16167
rect 6745 16133 6779 16167
rect 10333 16133 10367 16167
rect 10977 16133 11011 16167
rect 14381 16133 14415 16167
rect 14581 16133 14615 16167
rect 15117 16133 15151 16167
rect 1501 16065 1535 16099
rect 2789 16065 2823 16099
rect 4721 16065 4755 16099
rect 5089 16065 5123 16099
rect 6377 16065 6411 16099
rect 7757 16065 7791 16099
rect 9873 16065 9907 16099
rect 10793 16065 10827 16099
rect 11069 16065 11103 16099
rect 11713 16065 11747 16099
rect 12909 16065 12943 16099
rect 13093 16065 13127 16099
rect 13185 16065 13219 16099
rect 13277 16065 13311 16099
rect 13461 16065 13495 16099
rect 14841 16065 14875 16099
rect 14933 16065 14967 16099
rect 15393 16065 15427 16099
rect 15820 16065 15854 16099
rect 16037 16065 16071 16099
rect 16221 16065 16255 16099
rect 16313 16065 16347 16099
rect 2605 15997 2639 16031
rect 4629 15997 4663 16031
rect 9597 15997 9631 16031
rect 9965 15997 9999 16031
rect 15301 15997 15335 16031
rect 10609 15929 10643 15963
rect 15117 15929 15151 15963
rect 2973 15861 3007 15895
rect 4445 15861 4479 15895
rect 6745 15861 6779 15895
rect 6929 15861 6963 15895
rect 7665 15861 7699 15895
rect 10333 15861 10367 15895
rect 10517 15861 10551 15895
rect 11621 15861 11655 15895
rect 14565 15861 14599 15895
rect 15945 15861 15979 15895
rect 6469 15657 6503 15691
rect 9505 15657 9539 15691
rect 9689 15657 9723 15691
rect 11989 15657 12023 15691
rect 16405 15657 16439 15691
rect 17877 15657 17911 15691
rect 4445 15589 4479 15623
rect 9413 15589 9447 15623
rect 17693 15589 17727 15623
rect 1777 15521 1811 15555
rect 2053 15521 2087 15555
rect 7941 15521 7975 15555
rect 8217 15521 8251 15555
rect 10241 15521 10275 15555
rect 10517 15521 10551 15555
rect 15485 15521 15519 15555
rect 1685 15453 1719 15487
rect 3985 15453 4019 15487
rect 4169 15453 4203 15487
rect 4261 15453 4295 15487
rect 4353 15453 4387 15487
rect 4721 15453 4755 15487
rect 4813 15453 4847 15487
rect 4905 15453 4939 15487
rect 5089 15453 5123 15487
rect 6101 15453 6135 15487
rect 6285 15453 6319 15487
rect 8585 15453 8619 15487
rect 8769 15453 8803 15487
rect 9229 15453 9263 15487
rect 12725 15453 12759 15487
rect 12909 15453 12943 15487
rect 13093 15453 13127 15487
rect 14933 15453 14967 15487
rect 15301 15453 15335 15487
rect 15577 15453 15611 15487
rect 15761 15453 15795 15487
rect 16313 15453 16347 15487
rect 16497 15453 16531 15487
rect 17233 15453 17267 15487
rect 5273 15385 5307 15419
rect 9045 15385 9079 15419
rect 9873 15385 9907 15419
rect 12817 15385 12851 15419
rect 17417 15385 17451 15419
rect 17845 15385 17879 15419
rect 18061 15385 18095 15419
rect 6101 15317 6135 15351
rect 8769 15317 8803 15351
rect 9663 15317 9697 15351
rect 12541 15317 12575 15351
rect 17601 15317 17635 15351
rect 1593 15113 1627 15147
rect 2789 15113 2823 15147
rect 3249 15113 3283 15147
rect 5365 15113 5399 15147
rect 9045 15113 9079 15147
rect 10885 15113 10919 15147
rect 13461 15113 13495 15147
rect 17601 15113 17635 15147
rect 17693 15113 17727 15147
rect 5825 15045 5859 15079
rect 6025 15045 6059 15079
rect 8769 15045 8803 15079
rect 12633 15045 12667 15079
rect 16037 15045 16071 15079
rect 16221 15045 16255 15079
rect 1409 14977 1443 15011
rect 2237 14977 2271 15011
rect 2881 14977 2915 15011
rect 3341 14977 3375 15011
rect 3525 14977 3559 15011
rect 3709 14977 3743 15011
rect 3893 14977 3927 15011
rect 4445 14977 4479 15011
rect 4537 14977 4571 15011
rect 4813 14977 4847 15011
rect 6377 14977 6411 15011
rect 9137 14977 9171 15011
rect 9597 14977 9631 15011
rect 11713 14977 11747 15011
rect 13001 14977 13035 15011
rect 13277 14977 13311 15011
rect 13553 14977 13587 15011
rect 15209 14977 15243 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 16957 14977 16991 15011
rect 17141 14977 17175 15011
rect 17233 14977 17267 15011
rect 17509 14977 17543 15011
rect 18153 14977 18187 15011
rect 18337 14977 18371 15011
rect 18429 14977 18463 15011
rect 1685 14909 1719 14943
rect 2513 14909 2547 14943
rect 2973 14909 3007 14943
rect 3617 14909 3651 14943
rect 4169 14909 4203 14943
rect 4353 14909 4387 14943
rect 4629 14909 4663 14943
rect 5089 14909 5123 14943
rect 6653 14909 6687 14943
rect 8401 14909 8435 14943
rect 11989 14909 12023 14943
rect 15577 14909 15611 14943
rect 17325 14909 17359 14943
rect 2053 14841 2087 14875
rect 6193 14841 6227 14875
rect 15485 14841 15519 14875
rect 17877 14841 17911 14875
rect 17969 14841 18003 14875
rect 2145 14773 2179 14807
rect 2329 14773 2363 14807
rect 3065 14773 3099 14807
rect 4077 14773 4111 14807
rect 4905 14773 4939 14807
rect 6009 14773 6043 14807
rect 8677 14773 8711 14807
rect 12449 14773 12483 14807
rect 12633 14773 12667 14807
rect 13185 14773 13219 14807
rect 15347 14773 15381 14807
rect 15853 14773 15887 14807
rect 16405 14773 16439 14807
rect 3985 14569 4019 14603
rect 4261 14569 4295 14603
rect 4813 14569 4847 14603
rect 5089 14569 5123 14603
rect 6009 14569 6043 14603
rect 6745 14569 6779 14603
rect 9965 14569 9999 14603
rect 11915 14569 11949 14603
rect 16497 14569 16531 14603
rect 16681 14569 16715 14603
rect 17141 14569 17175 14603
rect 17325 14569 17359 14603
rect 17601 14569 17635 14603
rect 17785 14569 17819 14603
rect 1593 14501 1627 14535
rect 2513 14501 2547 14535
rect 2237 14433 2271 14467
rect 2697 14433 2731 14467
rect 4445 14433 4479 14467
rect 12173 14433 12207 14467
rect 15209 14433 15243 14467
rect 15945 14433 15979 14467
rect 16405 14433 16439 14467
rect 1409 14365 1443 14399
rect 3801 14365 3835 14399
rect 3985 14365 4019 14399
rect 4077 14365 4111 14399
rect 4261 14365 4295 14399
rect 4537 14365 4571 14399
rect 4905 14365 4939 14399
rect 6193 14365 6227 14399
rect 6377 14365 6411 14399
rect 13185 14365 13219 14399
rect 13553 14365 13587 14399
rect 13829 14365 13863 14399
rect 15853 14365 15887 14399
rect 16221 14365 16255 14399
rect 17049 14365 17083 14399
rect 18245 14365 18279 14399
rect 18521 14365 18555 14399
rect 8217 14297 8251 14331
rect 10149 14297 10183 14331
rect 10333 14297 10367 14331
rect 13277 14297 13311 14331
rect 13369 14297 13403 14331
rect 13737 14297 13771 14331
rect 17309 14297 17343 14331
rect 17509 14297 17543 14331
rect 17769 14297 17803 14331
rect 17969 14297 18003 14331
rect 10425 14229 10459 14263
rect 13001 14229 13035 14263
rect 16681 14229 16715 14263
rect 18061 14229 18095 14263
rect 18337 14229 18371 14263
rect 5825 14025 5859 14059
rect 7573 14025 7607 14059
rect 10175 14025 10209 14059
rect 10609 14025 10643 14059
rect 10701 14025 10735 14059
rect 12350 14025 12384 14059
rect 12909 14025 12943 14059
rect 15485 14025 15519 14059
rect 17049 14025 17083 14059
rect 18061 14025 18095 14059
rect 18429 14025 18463 14059
rect 6469 13957 6503 13991
rect 8953 13957 8987 13991
rect 9153 13957 9187 13991
rect 9965 13957 9999 13991
rect 10977 13957 11011 13991
rect 12449 13957 12483 13991
rect 13093 13957 13127 13991
rect 14013 13957 14047 13991
rect 15761 13957 15795 13991
rect 15853 13957 15887 13991
rect 16865 13957 16899 13991
rect 2053 13889 2087 13923
rect 2237 13889 2271 13923
rect 5733 13889 5767 13923
rect 6009 13889 6043 13923
rect 7665 13889 7699 13923
rect 10793 13889 10827 13923
rect 12173 13889 12207 13923
rect 12265 13889 12299 13923
rect 12725 13889 12759 13923
rect 12817 13889 12851 13923
rect 13369 13889 13403 13923
rect 13461 13889 13495 13923
rect 13921 13889 13955 13923
rect 15117 13889 15151 13923
rect 15301 13889 15335 13923
rect 15577 13889 15611 13923
rect 15945 13889 15979 13923
rect 16681 13889 16715 13923
rect 17601 13889 17635 13923
rect 17693 13889 17727 13923
rect 18153 13889 18187 13923
rect 12541 13821 12575 13855
rect 13737 13821 13771 13855
rect 13829 13821 13863 13855
rect 17785 13821 17819 13855
rect 18429 13821 18463 13855
rect 13185 13753 13219 13787
rect 16129 13753 16163 13787
rect 18245 13753 18279 13787
rect 2145 13685 2179 13719
rect 6193 13685 6227 13719
rect 9137 13685 9171 13719
rect 9321 13685 9355 13719
rect 10149 13685 10183 13719
rect 10333 13685 10367 13719
rect 10425 13685 10459 13719
rect 17509 13685 17543 13719
rect 17877 13685 17911 13719
rect 4445 13481 4479 13515
rect 5733 13481 5767 13515
rect 6377 13481 6411 13515
rect 8401 13481 8435 13515
rect 8677 13481 8711 13515
rect 10701 13481 10735 13515
rect 13277 13481 13311 13515
rect 13737 13481 13771 13515
rect 17141 13481 17175 13515
rect 2605 13413 2639 13447
rect 13001 13413 13035 13447
rect 2789 13345 2823 13379
rect 6653 13345 6687 13379
rect 8953 13345 8987 13379
rect 10885 13345 10919 13379
rect 17325 13345 17359 13379
rect 1409 13277 1443 13311
rect 1961 13277 1995 13311
rect 2145 13277 2179 13311
rect 3065 13277 3099 13311
rect 3341 13277 3375 13311
rect 3433 13277 3467 13311
rect 3893 13277 3927 13311
rect 4261 13277 4295 13311
rect 6009 13277 6043 13311
rect 8585 13277 8619 13311
rect 8769 13277 8803 13311
rect 12725 13277 12759 13311
rect 13001 13277 13035 13311
rect 13185 13277 13219 13311
rect 13461 13277 13495 13311
rect 13553 13277 13587 13311
rect 13829 13277 13863 13311
rect 17417 13277 17451 13311
rect 18521 13277 18555 13311
rect 2329 13209 2363 13243
rect 3249 13209 3283 13243
rect 4077 13209 4111 13243
rect 4169 13209 4203 13243
rect 5549 13209 5583 13243
rect 5749 13209 5783 13243
rect 6929 13209 6963 13243
rect 9229 13209 9263 13243
rect 11161 13209 11195 13243
rect 1593 13141 1627 13175
rect 2053 13141 2087 13175
rect 3617 13141 3651 13175
rect 5917 13141 5951 13175
rect 6377 13141 6411 13175
rect 6561 13141 6595 13175
rect 12633 13141 12667 13175
rect 18337 13141 18371 13175
rect 2421 12937 2455 12971
rect 4629 12937 4663 12971
rect 5641 12937 5675 12971
rect 5825 12937 5859 12971
rect 7849 12937 7883 12971
rect 9229 12937 9263 12971
rect 9781 12937 9815 12971
rect 10885 12937 10919 12971
rect 11805 12937 11839 12971
rect 14105 12937 14139 12971
rect 16129 12937 16163 12971
rect 18061 12937 18095 12971
rect 6745 12869 6779 12903
rect 7021 12869 7055 12903
rect 9597 12869 9631 12903
rect 10701 12869 10735 12903
rect 14222 12869 14256 12903
rect 18337 12869 18371 12903
rect 1593 12801 1627 12835
rect 2053 12801 2087 12835
rect 2513 12801 2547 12835
rect 3341 12801 3375 12835
rect 3801 12801 3835 12835
rect 3985 12801 4019 12835
rect 4077 12801 4111 12835
rect 4169 12801 4203 12835
rect 4353 12801 4387 12835
rect 4813 12801 4847 12835
rect 5089 12801 5123 12835
rect 5181 12801 5215 12835
rect 5365 12801 5399 12835
rect 5733 12801 5767 12835
rect 7205 12801 7239 12835
rect 7941 12801 7975 12835
rect 9413 12801 9447 12835
rect 9689 12801 9723 12835
rect 10333 12801 10367 12835
rect 11713 12801 11747 12835
rect 13737 12801 13771 12835
rect 15485 12801 15519 12835
rect 16313 12801 16347 12835
rect 16957 12801 16991 12835
rect 17417 12801 17451 12835
rect 18429 12801 18463 12835
rect 2145 12733 2179 12767
rect 2881 12733 2915 12767
rect 3433 12733 3467 12767
rect 4537 12733 4571 12767
rect 4997 12733 5031 12767
rect 5457 12733 5491 12767
rect 14013 12733 14047 12767
rect 15025 12733 15059 12767
rect 16497 12733 16531 12767
rect 16681 12733 16715 12767
rect 16865 12733 16899 12767
rect 17049 12733 17083 12767
rect 17141 12733 17175 12767
rect 17785 12733 17819 12767
rect 2789 12665 2823 12699
rect 6377 12665 6411 12699
rect 7389 12665 7423 12699
rect 14381 12665 14415 12699
rect 14473 12665 14507 12699
rect 14841 12665 14875 12699
rect 14933 12665 14967 12699
rect 1685 12597 1719 12631
rect 2651 12597 2685 12631
rect 2973 12597 3007 12631
rect 6009 12597 6043 12631
rect 6745 12597 6779 12631
rect 6929 12597 6963 12631
rect 10701 12597 10735 12631
rect 15117 12597 15151 12631
rect 15577 12597 15611 12631
rect 17582 12597 17616 12631
rect 17693 12597 17727 12631
rect 1593 12393 1627 12427
rect 3617 12393 3651 12427
rect 5089 12393 5123 12427
rect 8217 12393 8251 12427
rect 10517 12393 10551 12427
rect 14473 12393 14507 12427
rect 16129 12393 16163 12427
rect 17509 12393 17543 12427
rect 2605 12325 2639 12359
rect 15117 12325 15151 12359
rect 18337 12325 18371 12359
rect 4169 12257 4203 12291
rect 4261 12257 4295 12291
rect 5457 12257 5491 12291
rect 10701 12257 10735 12291
rect 14657 12257 14691 12291
rect 14749 12257 14783 12291
rect 14933 12257 14967 12291
rect 15577 12257 15611 12291
rect 1409 12189 1443 12223
rect 2145 12189 2179 12223
rect 2421 12189 2455 12223
rect 2697 12189 2731 12223
rect 2881 12189 2915 12223
rect 3433 12189 3467 12223
rect 3893 12189 3927 12223
rect 4077 12189 4111 12223
rect 4445 12189 4479 12223
rect 4721 12189 4755 12223
rect 4905 12189 4939 12223
rect 5181 12189 5215 12223
rect 5273 12189 5307 12223
rect 6469 12189 6503 12223
rect 8493 12189 8527 12223
rect 10057 12189 10091 12223
rect 10149 12189 10183 12223
rect 10333 12189 10367 12223
rect 11253 12189 11287 12223
rect 11805 12189 11839 12223
rect 14841 12189 14875 12223
rect 15485 12189 15519 12223
rect 15761 12189 15795 12223
rect 15945 12189 15979 12223
rect 16037 12189 16071 12223
rect 17601 12189 17635 12223
rect 18521 12189 18555 12223
rect 3249 12121 3283 12155
rect 4629 12121 4663 12155
rect 6745 12121 6779 12155
rect 8401 12121 8435 12155
rect 2237 12053 2271 12087
rect 3065 12053 3099 12087
rect 5457 12053 5491 12087
rect 11897 12053 11931 12087
rect 15761 12053 15795 12087
rect 1593 11849 1627 11883
rect 7573 11849 7607 11883
rect 8033 11781 8067 11815
rect 9597 11781 9631 11815
rect 10793 11781 10827 11815
rect 1409 11713 1443 11747
rect 2237 11713 2271 11747
rect 3985 11713 4019 11747
rect 4078 11713 4112 11747
rect 9873 11713 9907 11747
rect 10057 11713 10091 11747
rect 11529 11713 11563 11747
rect 13553 11713 13587 11747
rect 13829 11713 13863 11747
rect 14013 11713 14047 11747
rect 14105 11713 14139 11747
rect 14289 11713 14323 11747
rect 15577 11713 15611 11747
rect 15761 11713 15795 11747
rect 15853 11713 15887 11747
rect 10425 11645 10459 11679
rect 11805 11645 11839 11679
rect 13369 11645 13403 11679
rect 13737 11645 13771 11679
rect 7389 11577 7423 11611
rect 7941 11577 7975 11611
rect 10977 11577 11011 11611
rect 2145 11509 2179 11543
rect 4169 11509 4203 11543
rect 7573 11509 7607 11543
rect 9965 11509 9999 11543
rect 10793 11509 10827 11543
rect 13277 11509 13311 11543
rect 13829 11509 13863 11543
rect 14105 11509 14139 11543
rect 15393 11509 15427 11543
rect 1409 11305 1443 11339
rect 4629 11305 4663 11339
rect 5549 11305 5583 11339
rect 8953 11305 8987 11339
rect 10793 11305 10827 11339
rect 11805 11305 11839 11339
rect 13921 11305 13955 11339
rect 16773 11305 16807 11339
rect 9229 11237 9263 11271
rect 16589 11237 16623 11271
rect 2881 11169 2915 11203
rect 3157 11169 3191 11203
rect 5825 11169 5859 11203
rect 7573 11169 7607 11203
rect 9321 11169 9355 11203
rect 9413 11169 9447 11203
rect 9689 11169 9723 11203
rect 10149 11169 10183 11203
rect 16221 11169 16255 11203
rect 16405 11169 16439 11203
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4169 11101 4203 11135
rect 4445 11101 4479 11135
rect 4599 11101 4633 11135
rect 5181 11101 5215 11135
rect 7941 11101 7975 11135
rect 9137 11101 9171 11135
rect 9597 11101 9631 11135
rect 9873 11101 9907 11135
rect 10057 11101 10091 11135
rect 10425 11101 10459 11135
rect 11069 11101 11103 11135
rect 11345 11101 11379 11135
rect 13185 11101 13219 11135
rect 13369 11101 13403 11135
rect 13461 11101 13495 11135
rect 13553 11101 13587 11135
rect 13737 11101 13771 11135
rect 16129 11101 16163 11135
rect 16313 11101 16347 11135
rect 17877 11101 17911 11135
rect 18245 11101 18279 11135
rect 18521 11101 18555 11135
rect 4077 11033 4111 11067
rect 5549 11033 5583 11067
rect 6101 11033 6135 11067
rect 7849 11033 7883 11067
rect 11437 11033 11471 11067
rect 11621 11033 11655 11067
rect 16757 11033 16791 11067
rect 16957 11033 16991 11067
rect 4353 10965 4387 10999
rect 5733 10965 5767 10999
rect 10609 10965 10643 10999
rect 10977 10965 11011 10999
rect 11161 10965 11195 10999
rect 15945 10965 15979 10999
rect 17785 10965 17819 10999
rect 18061 10965 18095 10999
rect 18337 10965 18371 10999
rect 1593 10761 1627 10795
rect 2789 10761 2823 10795
rect 5549 10761 5583 10795
rect 9229 10761 9263 10795
rect 11161 10761 11195 10795
rect 13001 10761 13035 10795
rect 13737 10761 13771 10795
rect 16865 10761 16899 10795
rect 5917 10693 5951 10727
rect 9689 10693 9723 10727
rect 10793 10693 10827 10727
rect 10993 10693 11027 10727
rect 12817 10693 12851 10727
rect 16313 10693 16347 10727
rect 1409 10625 1443 10659
rect 2421 10625 2455 10659
rect 3985 10625 4019 10659
rect 4169 10625 4203 10659
rect 4445 10625 4479 10659
rect 5273 10625 5307 10659
rect 5733 10625 5767 10659
rect 8769 10625 8803 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 10057 10625 10091 10659
rect 10425 10625 10459 10659
rect 10609 10625 10643 10659
rect 10701 10625 10735 10659
rect 12173 10625 12207 10659
rect 12357 10625 12391 10659
rect 12633 10625 12667 10659
rect 13645 10625 13679 10659
rect 13921 10625 13955 10659
rect 14013 10625 14047 10659
rect 14289 10625 14323 10659
rect 15117 10625 15151 10659
rect 15301 10625 15335 10659
rect 15485 10625 15519 10659
rect 15853 10625 15887 10659
rect 16129 10625 16163 10659
rect 16405 10625 16439 10659
rect 17049 10625 17083 10659
rect 17877 10625 17911 10659
rect 18337 10625 18371 10659
rect 2513 10557 2547 10591
rect 5089 10557 5123 10591
rect 6377 10557 6411 10591
rect 6653 10557 6687 10591
rect 13369 10557 13403 10591
rect 15577 10557 15611 10591
rect 15945 10557 15979 10591
rect 17141 10557 17175 10591
rect 17233 10557 17267 10591
rect 17325 10557 17359 10591
rect 17785 10557 17819 10591
rect 8861 10489 8895 10523
rect 12541 10489 12575 10523
rect 14197 10489 14231 10523
rect 15761 10489 15795 10523
rect 17509 10489 17543 10523
rect 4629 10421 4663 10455
rect 5457 10421 5491 10455
rect 8125 10421 8159 10455
rect 9505 10421 9539 10455
rect 9689 10421 9723 10455
rect 10241 10421 10275 10455
rect 10977 10421 11011 10455
rect 13093 10421 13127 10455
rect 13553 10421 13587 10455
rect 15209 10421 15243 10455
rect 15485 10421 15519 10455
rect 18245 10421 18279 10455
rect 2697 10217 2731 10251
rect 9045 10217 9079 10251
rect 9762 10217 9796 10251
rect 11253 10217 11287 10251
rect 12909 10217 12943 10251
rect 13369 10217 13403 10251
rect 15025 10217 15059 10251
rect 16221 10217 16255 10251
rect 16313 10217 16347 10251
rect 16865 10217 16899 10251
rect 17969 10217 18003 10251
rect 5457 10149 5491 10183
rect 13185 10149 13219 10183
rect 15209 10149 15243 10183
rect 17509 10149 17543 10183
rect 18245 10149 18279 10183
rect 2513 10081 2547 10115
rect 9505 10081 9539 10115
rect 12817 10081 12851 10115
rect 14565 10081 14599 10115
rect 15117 10081 15151 10115
rect 15338 10081 15372 10115
rect 17785 10081 17819 10115
rect 1409 10013 1443 10047
rect 2789 10013 2823 10047
rect 4721 10013 4755 10047
rect 5089 10013 5123 10047
rect 5273 10013 5307 10047
rect 5917 10013 5951 10047
rect 6561 10013 6595 10047
rect 8033 10013 8067 10047
rect 8677 10013 8711 10047
rect 9137 10013 9171 10047
rect 11529 10013 11563 10047
rect 13001 10013 13035 10047
rect 13093 10013 13127 10047
rect 13369 10013 13403 10047
rect 13553 10013 13587 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14657 10013 14691 10047
rect 15577 10013 15611 10047
rect 15761 10013 15795 10047
rect 15853 10013 15887 10047
rect 15945 10013 15979 10047
rect 16313 10013 16347 10047
rect 16405 10013 16439 10047
rect 17049 10013 17083 10047
rect 17325 10013 17359 10047
rect 18061 10013 18095 10047
rect 18337 10013 18371 10047
rect 6653 9945 6687 9979
rect 6837 9945 6871 9979
rect 7481 9945 7515 9979
rect 8401 9945 8435 9979
rect 11437 9945 11471 9979
rect 13829 9945 13863 9979
rect 14105 9945 14139 9979
rect 15485 9945 15519 9979
rect 1593 9877 1627 9911
rect 2053 9877 2087 9911
rect 4261 9877 4295 9911
rect 5273 9877 5307 9911
rect 6101 9877 6135 9911
rect 7021 9877 7055 9911
rect 16681 9877 16715 9911
rect 17233 9877 17267 9911
rect 6193 9673 6227 9707
rect 10333 9673 10367 9707
rect 13645 9673 13679 9707
rect 15209 9673 15243 9707
rect 15853 9673 15887 9707
rect 18337 9673 18371 9707
rect 1777 9605 1811 9639
rect 2697 9605 2731 9639
rect 3275 9605 3309 9639
rect 5825 9605 5859 9639
rect 6041 9605 6075 9639
rect 10425 9605 10459 9639
rect 10625 9605 10659 9639
rect 11069 9605 11103 9639
rect 13553 9605 13587 9639
rect 15577 9605 15611 9639
rect 18245 9605 18279 9639
rect 1501 9537 1535 9571
rect 1593 9537 1627 9571
rect 1869 9537 1903 9571
rect 1961 9537 1995 9571
rect 2513 9537 2547 9571
rect 3400 9537 3434 9571
rect 3617 9537 3651 9571
rect 3801 9537 3835 9571
rect 4169 9537 4203 9571
rect 10149 9537 10183 9571
rect 10333 9537 10367 9571
rect 11253 9537 11287 9571
rect 13829 9537 13863 9571
rect 13921 9537 13955 9571
rect 14013 9537 14047 9571
rect 14197 9537 14231 9571
rect 14933 9537 14967 9571
rect 15301 9537 15335 9571
rect 15485 9537 15519 9571
rect 15674 9537 15708 9571
rect 16221 9537 16255 9571
rect 17969 9537 18003 9571
rect 18521 9537 18555 9571
rect 1777 9469 1811 9503
rect 2329 9469 2363 9503
rect 2881 9469 2915 9503
rect 3893 9469 3927 9503
rect 3985 9469 4019 9503
rect 11529 9469 11563 9503
rect 11805 9469 11839 9503
rect 15209 9469 15243 9503
rect 15393 9469 15427 9503
rect 16129 9469 16163 9503
rect 18061 9469 18095 9503
rect 2237 9401 2271 9435
rect 3525 9401 3559 9435
rect 10885 9401 10919 9435
rect 15025 9401 15059 9435
rect 17785 9401 17819 9435
rect 1869 9333 1903 9367
rect 2973 9333 3007 9367
rect 4353 9333 4387 9367
rect 6009 9333 6043 9367
rect 10609 9333 10643 9367
rect 10793 9333 10827 9367
rect 16221 9333 16255 9367
rect 18245 9333 18279 9367
rect 1593 9129 1627 9163
rect 3065 9129 3099 9163
rect 4905 9129 4939 9163
rect 8953 9129 8987 9163
rect 11989 9129 12023 9163
rect 16773 9129 16807 9163
rect 17877 9129 17911 9163
rect 17969 9129 18003 9163
rect 18429 9129 18463 9163
rect 2513 9061 2547 9095
rect 4721 9061 4755 9095
rect 5733 9061 5767 9095
rect 8309 9061 8343 9095
rect 8677 9061 8711 9095
rect 2237 8993 2271 9027
rect 2881 8993 2915 9027
rect 3617 8993 3651 9027
rect 4077 8993 4111 9027
rect 4169 8993 4203 9027
rect 5825 8993 5859 9027
rect 8401 8993 8435 9027
rect 10701 8993 10735 9027
rect 17233 8993 17267 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 1777 8925 1811 8959
rect 2145 8925 2179 8959
rect 2789 8925 2823 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 3985 8925 4019 8959
rect 4261 8925 4295 8959
rect 5181 8925 5215 8959
rect 5365 8925 5399 8959
rect 6009 8925 6043 8959
rect 6193 8925 6227 8959
rect 7113 8925 7147 8959
rect 7206 8925 7240 8959
rect 7389 8925 7423 8959
rect 7578 8925 7612 8959
rect 8180 8925 8214 8959
rect 9137 8925 9171 8959
rect 9321 8925 9355 8959
rect 9413 8925 9447 8959
rect 10425 8925 10459 8959
rect 11897 8925 11931 8959
rect 16773 8925 16807 8959
rect 16957 8925 16991 8959
rect 18153 8925 18187 8959
rect 18245 8925 18279 8959
rect 3065 8857 3099 8891
rect 5089 8857 5123 8891
rect 5457 8857 5491 8891
rect 7481 8857 7515 8891
rect 8033 8857 8067 8891
rect 17718 8857 17752 8891
rect 18429 8857 18463 8891
rect 2605 8789 2639 8823
rect 3801 8789 3835 8823
rect 4889 8789 4923 8823
rect 5549 8789 5583 8823
rect 7757 8789 7791 8823
rect 17509 8789 17543 8823
rect 17601 8789 17635 8823
rect 4353 8585 4387 8619
rect 4997 8585 5031 8619
rect 8309 8585 8343 8619
rect 9321 8585 9355 8619
rect 10609 8585 10643 8619
rect 13277 8585 13311 8619
rect 14473 8585 14507 8619
rect 16865 8585 16899 8619
rect 17785 8585 17819 8619
rect 3985 8517 4019 8551
rect 4077 8517 4111 8551
rect 7481 8517 7515 8551
rect 8953 8517 8987 8551
rect 9137 8517 9171 8551
rect 10057 8517 10091 8551
rect 11989 8517 12023 8551
rect 18429 8517 18463 8551
rect 2329 8449 2363 8483
rect 3525 8449 3559 8483
rect 3801 8449 3835 8483
rect 4169 8449 4203 8483
rect 4721 8449 4755 8483
rect 4813 8449 4847 8483
rect 5733 8449 5767 8483
rect 5917 8449 5951 8483
rect 6009 8449 6043 8483
rect 6469 8449 6503 8483
rect 6745 8449 6779 8483
rect 6929 8449 6963 8483
rect 7021 8449 7055 8483
rect 7297 8449 7331 8483
rect 7941 8449 7975 8483
rect 8125 8449 8159 8483
rect 8806 8449 8840 8483
rect 9045 8449 9079 8483
rect 9229 8449 9263 8483
rect 9505 8449 9539 8483
rect 9597 8449 9631 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 10517 8449 10551 8483
rect 10701 8449 10735 8483
rect 11805 8449 11839 8483
rect 13552 8449 13586 8483
rect 13645 8449 13679 8483
rect 13737 8449 13771 8483
rect 13921 8449 13955 8483
rect 14289 8449 14323 8483
rect 17141 8449 17175 8483
rect 17325 8449 17359 8483
rect 17601 8449 17635 8483
rect 17693 8449 17727 8483
rect 17871 8449 17905 8483
rect 17969 8449 18003 8483
rect 1409 8381 1443 8415
rect 1685 8381 1719 8415
rect 2697 8381 2731 8415
rect 3433 8381 3467 8415
rect 4537 8381 4571 8415
rect 4629 8381 4663 8415
rect 6101 8381 6135 8415
rect 7113 8381 7147 8415
rect 8585 8381 8619 8415
rect 14013 8381 14047 8415
rect 14105 8381 14139 8415
rect 2494 8313 2528 8347
rect 3157 8313 3191 8347
rect 6561 8313 6595 8347
rect 8033 8313 8067 8347
rect 17233 8313 17267 8347
rect 2605 8245 2639 8279
rect 2973 8245 3007 8279
rect 3341 8245 3375 8279
rect 5825 8245 5859 8279
rect 8677 8245 8711 8279
rect 11621 8245 11655 8279
rect 17417 8245 17451 8279
rect 18061 8245 18095 8279
rect 18337 8245 18371 8279
rect 2881 8041 2915 8075
rect 4537 8041 4571 8075
rect 7573 8041 7607 8075
rect 8493 8041 8527 8075
rect 9229 8041 9263 8075
rect 10149 8041 10183 8075
rect 10977 8041 11011 8075
rect 14197 8041 14231 8075
rect 14565 8041 14599 8075
rect 15577 8041 15611 8075
rect 18337 8041 18371 8075
rect 7297 7973 7331 8007
rect 14657 7973 14691 8007
rect 15025 7973 15059 8007
rect 15117 7973 15151 8007
rect 17325 7973 17359 8007
rect 17509 7973 17543 8007
rect 2605 7905 2639 7939
rect 3157 7905 3191 7939
rect 4629 7905 4663 7939
rect 5089 7905 5123 7939
rect 6745 7905 6779 7939
rect 11253 7905 11287 7939
rect 13461 7905 13495 7939
rect 13553 7905 13587 7939
rect 16681 7905 16715 7939
rect 1409 7837 1443 7871
rect 1685 7837 1719 7871
rect 2513 7837 2547 7871
rect 3341 7837 3375 7871
rect 3985 7837 4019 7871
rect 4169 7837 4203 7871
rect 4353 7837 4387 7871
rect 4813 7837 4847 7871
rect 4905 7837 4939 7871
rect 5181 7837 5215 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 6193 7837 6227 7871
rect 6377 7837 6411 7871
rect 7711 7837 7745 7871
rect 7941 7837 7975 7871
rect 8069 7837 8103 7871
rect 8217 7837 8251 7871
rect 8309 7837 8343 7871
rect 8402 7837 8436 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 9505 7837 9539 7871
rect 9597 7837 9631 7871
rect 10024 7837 10058 7871
rect 10241 7837 10275 7871
rect 10609 7837 10643 7871
rect 14473 7837 14507 7871
rect 14933 7837 14967 7871
rect 15577 7837 15611 7871
rect 15761 7837 15795 7871
rect 16037 7837 16071 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 17141 7837 17175 7871
rect 17417 7837 17451 7871
rect 18061 7837 18095 7871
rect 18429 7837 18463 7871
rect 4261 7769 4295 7803
rect 7021 7769 7055 7803
rect 7849 7769 7883 7803
rect 10333 7769 10367 7803
rect 11529 7769 11563 7803
rect 15485 7769 15519 7803
rect 15945 7769 15979 7803
rect 17693 7769 17727 7803
rect 17877 7769 17911 7803
rect 3525 7701 3559 7735
rect 7481 7701 7515 7735
rect 9045 7701 9079 7735
rect 9965 7701 9999 7735
rect 10977 7701 11011 7735
rect 11161 7701 11195 7735
rect 13001 7701 13035 7735
rect 13277 7701 13311 7735
rect 13921 7701 13955 7735
rect 14841 7701 14875 7735
rect 16221 7701 16255 7735
rect 16589 7701 16623 7735
rect 2881 7497 2915 7531
rect 5273 7497 5307 7531
rect 6653 7497 6687 7531
rect 9413 7497 9447 7531
rect 10885 7497 10919 7531
rect 11621 7497 11655 7531
rect 12357 7497 12391 7531
rect 13461 7497 13495 7531
rect 13921 7497 13955 7531
rect 18337 7497 18371 7531
rect 9597 7429 9631 7463
rect 11897 7429 11931 7463
rect 15301 7429 15335 7463
rect 17509 7429 17543 7463
rect 18153 7429 18187 7463
rect 2605 7361 2639 7395
rect 4905 7361 4939 7395
rect 6928 7361 6962 7395
rect 7021 7361 7055 7395
rect 7113 7361 7147 7395
rect 9321 7361 9355 7395
rect 11805 7361 11839 7395
rect 11989 7361 12023 7395
rect 12265 7361 12299 7395
rect 13736 7361 13770 7395
rect 13829 7361 13863 7395
rect 14105 7361 14139 7395
rect 14289 7361 14323 7395
rect 14381 7361 14415 7395
rect 14565 7361 14599 7395
rect 14841 7361 14875 7395
rect 14933 7361 14967 7395
rect 15209 7361 15243 7395
rect 15485 7361 15519 7395
rect 16129 7361 16163 7395
rect 16497 7361 16531 7395
rect 16681 7361 16715 7395
rect 16773 7361 16807 7395
rect 17969 7361 18003 7395
rect 2881 7293 2915 7327
rect 12173 7293 12207 7327
rect 15669 7293 15703 7327
rect 16037 7293 16071 7327
rect 2697 7225 2731 7259
rect 14197 7225 14231 7259
rect 14657 7225 14691 7259
rect 16313 7225 16347 7259
rect 17877 7225 17911 7259
rect 5273 7157 5307 7191
rect 5457 7157 5491 7191
rect 15117 7157 15151 7191
rect 16957 7157 16991 7191
rect 17325 7157 17359 7191
rect 17509 7157 17543 7191
rect 5076 6953 5110 6987
rect 6561 6953 6595 6987
rect 12081 6953 12115 6987
rect 12265 6953 12299 6987
rect 17049 6953 17083 6987
rect 11391 6885 11425 6919
rect 11529 6885 11563 6919
rect 16957 6885 16991 6919
rect 4813 6817 4847 6851
rect 7113 6817 7147 6851
rect 11621 6817 11655 6851
rect 6837 6749 6871 6783
rect 9321 6749 9355 6783
rect 9873 6749 9907 6783
rect 10149 6749 10183 6783
rect 10425 6749 10459 6783
rect 10885 6749 10919 6783
rect 11989 6749 12023 6783
rect 13177 6743 13211 6777
rect 16681 6749 16715 6783
rect 17233 6749 17267 6783
rect 17693 6749 17727 6783
rect 18153 6749 18187 6783
rect 4537 6681 4571 6715
rect 4721 6681 4755 6715
rect 6745 6681 6779 6715
rect 8769 6681 8803 6715
rect 11253 6681 11287 6715
rect 12449 6681 12483 6715
rect 16773 6681 16807 6715
rect 16957 6681 16991 6715
rect 4353 6613 4387 6647
rect 9505 6613 9539 6647
rect 11069 6613 11103 6647
rect 12239 6613 12273 6647
rect 13277 6613 13311 6647
rect 17325 6613 17359 6647
rect 6193 6409 6227 6443
rect 7573 6409 7607 6443
rect 10517 6409 10551 6443
rect 12081 6409 12115 6443
rect 13921 6409 13955 6443
rect 16405 6409 16439 6443
rect 17049 6409 17083 6443
rect 6469 6341 6503 6375
rect 7113 6341 7147 6375
rect 9229 6341 9263 6375
rect 10333 6341 10367 6375
rect 11897 6341 11931 6375
rect 12449 6341 12483 6375
rect 15209 6341 15243 6375
rect 4445 6273 4479 6307
rect 6561 6273 6595 6307
rect 6837 6273 6871 6307
rect 7297 6273 7331 6307
rect 7757 6273 7791 6307
rect 8217 6273 8251 6307
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 8861 6273 8895 6307
rect 9137 6273 9171 6307
rect 9873 6273 9907 6307
rect 10057 6273 10091 6307
rect 10149 6273 10183 6307
rect 10425 6273 10459 6307
rect 10701 6273 10735 6307
rect 10977 6273 11011 6307
rect 11161 6273 11195 6307
rect 11529 6273 11563 6307
rect 15025 6273 15059 6307
rect 15301 6273 15335 6307
rect 15393 6273 15427 6307
rect 15853 6273 15887 6307
rect 15945 6273 15979 6307
rect 16221 6273 16255 6307
rect 16313 6273 16347 6307
rect 16497 6273 16531 6307
rect 17417 6273 17451 6307
rect 18245 6273 18279 6307
rect 4721 6205 4755 6239
rect 6929 6205 6963 6239
rect 7941 6205 7975 6239
rect 9045 6205 9079 6239
rect 12173 6205 12207 6239
rect 17325 6205 17359 6239
rect 18521 6205 18555 6239
rect 8033 6137 8067 6171
rect 9965 6137 9999 6171
rect 16129 6137 16163 6171
rect 7481 6069 7515 6103
rect 8493 6069 8527 6103
rect 10885 6069 10919 6103
rect 10977 6069 11011 6103
rect 11897 6069 11931 6103
rect 15577 6069 15611 6103
rect 15669 6069 15703 6103
rect 4721 5865 4755 5899
rect 10333 5865 10367 5899
rect 11989 5865 12023 5899
rect 15117 5865 15151 5899
rect 15301 5865 15335 5899
rect 18337 5865 18371 5899
rect 4537 5797 4571 5831
rect 5089 5797 5123 5831
rect 8401 5797 8435 5831
rect 11161 5797 11195 5831
rect 15393 5797 15427 5831
rect 15853 5797 15887 5831
rect 7665 5729 7699 5763
rect 9689 5729 9723 5763
rect 10057 5729 10091 5763
rect 10977 5729 11011 5763
rect 14657 5729 14691 5763
rect 15209 5729 15243 5763
rect 15761 5729 15795 5763
rect 7297 5661 7331 5695
rect 7481 5661 7515 5695
rect 7849 5661 7883 5695
rect 8125 5661 8159 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 9321 5661 9355 5695
rect 9505 5661 9539 5695
rect 9597 5661 9631 5695
rect 9873 5661 9907 5695
rect 10241 5661 10275 5695
rect 10517 5661 10551 5695
rect 10793 5661 10827 5695
rect 11161 5661 11195 5695
rect 12173 5661 12207 5695
rect 12633 5661 12667 5695
rect 12725 5661 12759 5695
rect 13553 5661 13587 5695
rect 14105 5661 14139 5695
rect 14565 5661 14599 5695
rect 14749 5661 14783 5695
rect 15991 5661 16025 5695
rect 16132 5661 16166 5695
rect 16404 5661 16438 5695
rect 16490 5661 16524 5695
rect 16589 5661 16623 5695
rect 16773 5661 16807 5695
rect 16957 5661 16991 5695
rect 18521 5661 18555 5695
rect 4721 5593 4755 5627
rect 7389 5593 7423 5627
rect 8033 5593 8067 5627
rect 8401 5593 8435 5627
rect 8585 5593 8619 5627
rect 10701 5593 10735 5627
rect 12357 5593 12391 5627
rect 12449 5593 12483 5627
rect 13001 5593 13035 5627
rect 14289 5593 14323 5627
rect 16221 5593 16255 5627
rect 16865 5593 16899 5627
rect 8217 5525 8251 5559
rect 10885 5525 10919 5559
rect 14473 5525 14507 5559
rect 17141 5525 17175 5559
rect 9229 5321 9263 5355
rect 10425 5321 10459 5355
rect 15577 5321 15611 5355
rect 16313 5321 16347 5355
rect 4813 5253 4847 5287
rect 8861 5253 8895 5287
rect 9965 5253 9999 5287
rect 12357 5253 12391 5287
rect 14657 5253 14691 5287
rect 4997 5185 5031 5219
rect 5273 5185 5307 5219
rect 5457 5185 5491 5219
rect 8217 5185 8251 5219
rect 8677 5185 8711 5219
rect 8953 5185 8987 5219
rect 9045 5185 9079 5219
rect 9689 5185 9723 5219
rect 9873 5185 9907 5219
rect 10057 5185 10091 5219
rect 10333 5185 10367 5219
rect 10517 5185 10551 5219
rect 11989 5185 12023 5219
rect 12633 5185 12667 5219
rect 14841 5185 14875 5219
rect 15025 5185 15059 5219
rect 15209 5185 15243 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 16129 5185 16163 5219
rect 8125 5117 8159 5151
rect 12909 5117 12943 5151
rect 14933 5117 14967 5151
rect 8585 5049 8619 5083
rect 10241 5049 10275 5083
rect 12541 5049 12575 5083
rect 15761 5049 15795 5083
rect 4629 4981 4663 5015
rect 5089 4981 5123 5015
rect 12357 4981 12391 5015
rect 15577 4981 15611 5015
rect 5917 4777 5951 4811
rect 9045 4777 9079 4811
rect 9505 4777 9539 4811
rect 13645 4777 13679 4811
rect 4169 4641 4203 4675
rect 6745 4573 6779 4607
rect 8953 4573 8987 4607
rect 9229 4573 9263 4607
rect 9321 4573 9355 4607
rect 12449 4573 12483 4607
rect 13553 4573 13587 4607
rect 4445 4505 4479 4539
rect 6653 4505 6687 4539
rect 6929 4505 6963 4539
rect 6377 4437 6411 4471
rect 6561 4437 6595 4471
rect 12357 4437 12391 4471
rect 4537 4233 4571 4267
rect 8309 4233 8343 4267
rect 11713 4233 11747 4267
rect 12081 4233 12115 4267
rect 4721 4165 4755 4199
rect 5549 4165 5583 4199
rect 5825 4165 5859 4199
rect 10517 4165 10551 4199
rect 11805 4165 11839 4199
rect 6055 4131 6089 4165
rect 5089 4097 5123 4131
rect 5365 4097 5399 4131
rect 6561 4097 6595 4131
rect 8493 4097 8527 4131
rect 8585 4097 8619 4131
rect 11529 4097 11563 4131
rect 11897 4097 11931 4131
rect 12173 4097 12207 4131
rect 12357 4097 12391 4131
rect 12449 4097 12483 4131
rect 12541 4097 12575 4131
rect 12909 4097 12943 4131
rect 6837 4029 6871 4063
rect 12817 4029 12851 4063
rect 13185 4029 13219 4063
rect 10149 3961 10183 3995
rect 10701 3961 10735 3995
rect 4721 3893 4755 3927
rect 5733 3893 5767 3927
rect 6009 3893 6043 3927
rect 6193 3893 6227 3927
rect 10517 3893 10551 3927
rect 14657 3893 14691 3927
rect 5181 3689 5215 3723
rect 6561 3689 6595 3723
rect 6745 3689 6779 3723
rect 8585 3689 8619 3723
rect 9505 3689 9539 3723
rect 9873 3689 9907 3723
rect 10057 3689 10091 3723
rect 12265 3689 12299 3723
rect 13829 3689 13863 3723
rect 6193 3621 6227 3655
rect 10425 3553 10459 3587
rect 11897 3553 11931 3587
rect 5273 3485 5307 3519
rect 6837 3485 6871 3519
rect 7021 3485 7055 3519
rect 9321 3485 9355 3519
rect 9413 3485 9447 3519
rect 9597 3485 9631 3519
rect 10149 3485 10183 3519
rect 12449 3485 12483 3519
rect 12633 3485 12667 3519
rect 12909 3485 12943 3519
rect 13093 3485 13127 3519
rect 13185 3485 13219 3519
rect 13737 3485 13771 3519
rect 6561 3417 6595 3451
rect 8401 3417 8435 3451
rect 8617 3417 8651 3451
rect 8953 3417 8987 3451
rect 9137 3417 9171 3451
rect 9689 3417 9723 3451
rect 9889 3417 9923 3451
rect 13369 3417 13403 3451
rect 7205 3349 7239 3383
rect 8769 3349 8803 3383
rect 12725 3349 12759 3383
rect 13553 3349 13587 3383
rect 14473 3145 14507 3179
rect 8861 3077 8895 3111
rect 10517 3077 10551 3111
rect 11621 3077 11655 3111
rect 12449 3077 12483 3111
rect 6745 3009 6779 3043
rect 8585 3009 8619 3043
rect 10701 3009 10735 3043
rect 10885 3009 10919 3043
rect 10977 3009 11011 3043
rect 11161 3009 11195 3043
rect 11253 3009 11287 3043
rect 11713 3009 11747 3043
rect 12081 3009 12115 3043
rect 12725 3009 12759 3043
rect 7021 2941 7055 2975
rect 8493 2941 8527 2975
rect 13001 2941 13035 2975
rect 10333 2873 10367 2907
rect 12633 2873 12667 2907
rect 12449 2805 12483 2839
rect 7021 2601 7055 2635
rect 7205 2601 7239 2635
rect 8033 2601 8067 2635
rect 8677 2601 8711 2635
rect 13737 2601 13771 2635
rect 6653 2533 6687 2567
rect 9413 2533 9447 2567
rect 10057 2465 10091 2499
rect 8125 2397 8159 2431
rect 8217 2397 8251 2431
rect 8493 2397 8527 2431
rect 9781 2397 9815 2431
rect 13645 2397 13679 2431
rect 7021 2329 7055 2363
rect 9229 2329 9263 2363
rect 8401 2261 8435 2295
<< metal1 >>
rect 14826 20680 14832 20732
rect 14884 20720 14890 20732
rect 16850 20720 16856 20732
rect 14884 20692 16856 20720
rect 14884 20680 14890 20692
rect 16850 20680 16856 20692
rect 16908 20680 16914 20732
rect 1104 19610 18860 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 18860 19610
rect 1104 19536 18860 19558
rect 14182 19456 14188 19508
rect 14240 19456 14246 19508
rect 15930 19456 15936 19508
rect 15988 19496 15994 19508
rect 16669 19499 16727 19505
rect 16669 19496 16681 19499
rect 15988 19468 16681 19496
rect 15988 19456 15994 19468
rect 16669 19465 16681 19468
rect 16715 19465 16727 19499
rect 16669 19459 16727 19465
rect 5629 19431 5687 19437
rect 5629 19397 5641 19431
rect 5675 19428 5687 19431
rect 5675 19400 6224 19428
rect 5675 19397 5687 19400
rect 5629 19391 5687 19397
rect 6196 19372 6224 19400
rect 7006 19388 7012 19440
rect 7064 19428 7070 19440
rect 7745 19431 7803 19437
rect 7745 19428 7757 19431
rect 7064 19400 7757 19428
rect 7064 19388 7070 19400
rect 7745 19397 7757 19400
rect 7791 19397 7803 19431
rect 14200 19428 14228 19456
rect 14200 19400 16528 19428
rect 7745 19391 7803 19397
rect 5905 19363 5963 19369
rect 5905 19360 5917 19363
rect 5736 19332 5917 19360
rect 5626 19184 5632 19236
rect 5684 19224 5690 19236
rect 5736 19224 5764 19332
rect 5905 19329 5917 19332
rect 5951 19329 5963 19363
rect 5905 19323 5963 19329
rect 6086 19320 6092 19372
rect 6144 19320 6150 19372
rect 6178 19320 6184 19372
rect 6236 19320 6242 19372
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 7377 19363 7435 19369
rect 7377 19360 7389 19363
rect 6512 19332 7389 19360
rect 6512 19320 6518 19332
rect 7377 19329 7389 19332
rect 7423 19329 7435 19363
rect 7377 19323 7435 19329
rect 11241 19363 11299 19369
rect 11241 19329 11253 19363
rect 11287 19360 11299 19363
rect 11330 19360 11336 19372
rect 11287 19332 11336 19360
rect 11287 19329 11299 19332
rect 11241 19323 11299 19329
rect 11330 19320 11336 19332
rect 11388 19320 11394 19372
rect 13262 19320 13268 19372
rect 13320 19320 13326 19372
rect 14182 19320 14188 19372
rect 14240 19320 14246 19372
rect 14277 19363 14335 19369
rect 14277 19329 14289 19363
rect 14323 19360 14335 19363
rect 15105 19363 15163 19369
rect 15105 19360 15117 19363
rect 14323 19332 15117 19360
rect 14323 19329 14335 19332
rect 14277 19323 14335 19329
rect 15105 19329 15117 19332
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15930 19320 15936 19372
rect 15988 19320 15994 19372
rect 16500 19369 16528 19400
rect 16209 19363 16267 19369
rect 16209 19329 16221 19363
rect 16255 19329 16267 19363
rect 16209 19323 16267 19329
rect 16485 19363 16543 19369
rect 16485 19329 16497 19363
rect 16531 19329 16543 19363
rect 16485 19323 16543 19329
rect 5810 19252 5816 19304
rect 5868 19292 5874 19304
rect 6365 19295 6423 19301
rect 6365 19292 6377 19295
rect 5868 19264 6377 19292
rect 5868 19252 5874 19264
rect 6365 19261 6377 19264
rect 6411 19261 6423 19295
rect 6365 19255 6423 19261
rect 6638 19252 6644 19304
rect 6696 19252 6702 19304
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12952 19264 13001 19292
rect 12952 19252 12958 19264
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 12989 19255 13047 19261
rect 14461 19295 14519 19301
rect 14461 19261 14473 19295
rect 14507 19261 14519 19295
rect 14461 19255 14519 19261
rect 9306 19224 9312 19236
rect 5684 19196 9312 19224
rect 5684 19184 5690 19196
rect 9306 19184 9312 19196
rect 9364 19184 9370 19236
rect 14274 19184 14280 19236
rect 14332 19224 14338 19236
rect 14476 19224 14504 19255
rect 15378 19252 15384 19304
rect 15436 19252 15442 19304
rect 15470 19252 15476 19304
rect 15528 19252 15534 19304
rect 16114 19224 16120 19236
rect 14332 19196 16120 19224
rect 14332 19184 14338 19196
rect 16114 19184 16120 19196
rect 16172 19184 16178 19236
rect 16224 19224 16252 19323
rect 16850 19320 16856 19372
rect 16908 19320 16914 19372
rect 16482 19224 16488 19236
rect 16224 19196 16488 19224
rect 11149 19159 11207 19165
rect 11149 19125 11161 19159
rect 11195 19156 11207 19159
rect 11238 19156 11244 19168
rect 11195 19128 11244 19156
rect 11195 19125 11207 19128
rect 11149 19119 11207 19125
rect 11238 19116 11244 19128
rect 11296 19116 11302 19168
rect 14366 19116 14372 19168
rect 14424 19116 14430 19168
rect 14826 19116 14832 19168
rect 14884 19156 14890 19168
rect 16224 19156 16252 19196
rect 16482 19184 16488 19196
rect 16540 19184 16546 19236
rect 14884 19128 16252 19156
rect 14884 19116 14890 19128
rect 16298 19116 16304 19168
rect 16356 19116 16362 19168
rect 1104 19066 18860 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 18860 19066
rect 1104 18992 18860 19014
rect 5810 18952 5816 18964
rect 4724 18924 5816 18952
rect 4614 18708 4620 18760
rect 4672 18708 4678 18760
rect 4724 18757 4752 18924
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 9858 18912 9864 18964
rect 9916 18952 9922 18964
rect 11330 18952 11336 18964
rect 9916 18924 11336 18952
rect 9916 18912 9922 18924
rect 11330 18912 11336 18924
rect 11388 18952 11394 18964
rect 11388 18924 11928 18952
rect 11388 18912 11394 18924
rect 5718 18776 5724 18828
rect 5776 18816 5782 18828
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 5776 18788 6837 18816
rect 5776 18776 5782 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 6825 18779 6883 18785
rect 9953 18819 10011 18825
rect 9953 18785 9965 18819
rect 9999 18816 10011 18819
rect 10778 18816 10784 18828
rect 9999 18788 10784 18816
rect 9999 18785 10011 18788
rect 9953 18779 10011 18785
rect 10778 18776 10784 18788
rect 10836 18816 10842 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 10836 18788 11805 18816
rect 10836 18776 10842 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11900 18816 11928 18924
rect 15378 18912 15384 18964
rect 15436 18952 15442 18964
rect 16485 18955 16543 18961
rect 16485 18952 16497 18955
rect 15436 18924 16497 18952
rect 15436 18912 15442 18924
rect 16114 18844 16120 18896
rect 16172 18844 16178 18896
rect 15930 18816 15936 18828
rect 11900 18788 13768 18816
rect 11793 18779 11851 18785
rect 4709 18751 4767 18757
rect 4709 18717 4721 18751
rect 4755 18717 4767 18751
rect 4709 18711 4767 18717
rect 5077 18751 5135 18757
rect 5077 18717 5089 18751
rect 5123 18717 5135 18751
rect 5077 18711 5135 18717
rect 4338 18640 4344 18692
rect 4396 18680 4402 18692
rect 5092 18680 5120 18711
rect 6454 18708 6460 18760
rect 6512 18708 6518 18760
rect 13740 18757 13768 18788
rect 15212 18788 15936 18816
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18717 13783 18751
rect 13725 18711 13783 18717
rect 14182 18708 14188 18760
rect 14240 18708 14246 18760
rect 14274 18708 14280 18760
rect 14332 18748 14338 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 14332 18720 14473 18748
rect 14332 18708 14338 18720
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 14461 18711 14519 18717
rect 14826 18708 14832 18760
rect 14884 18708 14890 18760
rect 4396 18652 5120 18680
rect 4396 18640 4402 18652
rect 4614 18572 4620 18624
rect 4672 18612 4678 18624
rect 4893 18615 4951 18621
rect 4893 18612 4905 18615
rect 4672 18584 4905 18612
rect 4672 18572 4678 18584
rect 4893 18581 4905 18584
rect 4939 18581 4951 18615
rect 5092 18612 5120 18652
rect 5258 18640 5264 18692
rect 5316 18680 5322 18692
rect 5353 18683 5411 18689
rect 5353 18680 5365 18683
rect 5316 18652 5365 18680
rect 5316 18640 5322 18652
rect 5353 18649 5365 18652
rect 5399 18649 5411 18683
rect 5353 18643 5411 18649
rect 10226 18640 10232 18692
rect 10284 18640 10290 18692
rect 11238 18640 11244 18692
rect 11296 18640 11302 18692
rect 12066 18640 12072 18692
rect 12124 18640 12130 18692
rect 13817 18683 13875 18689
rect 13817 18680 13829 18683
rect 13294 18652 13829 18680
rect 13817 18649 13829 18652
rect 13863 18649 13875 18683
rect 14200 18680 14228 18708
rect 15212 18680 15240 18788
rect 15930 18776 15936 18788
rect 15988 18816 15994 18828
rect 16025 18819 16083 18825
rect 16025 18816 16037 18819
rect 15988 18788 16037 18816
rect 15988 18776 15994 18788
rect 16025 18785 16037 18788
rect 16071 18785 16083 18819
rect 16025 18779 16083 18785
rect 16298 18757 16304 18760
rect 15381 18751 15439 18757
rect 15381 18717 15393 18751
rect 15427 18748 15439 18751
rect 16246 18751 16304 18757
rect 16246 18748 16258 18751
rect 15427 18720 16258 18748
rect 15427 18717 15439 18720
rect 15381 18711 15439 18717
rect 16246 18717 16258 18720
rect 16292 18717 16304 18751
rect 16246 18711 16304 18717
rect 14200 18652 15240 18680
rect 13817 18643 13875 18649
rect 15286 18640 15292 18692
rect 15344 18640 15350 18692
rect 6730 18612 6736 18624
rect 5092 18584 6736 18612
rect 4893 18575 4951 18581
rect 6730 18572 6736 18584
rect 6788 18572 6794 18624
rect 11698 18572 11704 18624
rect 11756 18572 11762 18624
rect 13078 18572 13084 18624
rect 13136 18612 13142 18624
rect 13538 18612 13544 18624
rect 13136 18584 13544 18612
rect 13136 18572 13142 18584
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 13722 18572 13728 18624
rect 13780 18612 13786 18624
rect 15396 18612 15424 18711
rect 16298 18708 16304 18711
rect 16356 18708 16362 18760
rect 16408 18757 16436 18924
rect 16485 18921 16497 18924
rect 16531 18921 16543 18955
rect 16485 18915 16543 18921
rect 16393 18751 16451 18757
rect 16393 18717 16405 18751
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 16482 18708 16488 18760
rect 16540 18748 16546 18760
rect 16669 18751 16727 18757
rect 16669 18748 16681 18751
rect 16540 18720 16681 18748
rect 16540 18708 16546 18720
rect 16669 18717 16681 18720
rect 16715 18717 16727 18751
rect 16669 18711 16727 18717
rect 13780 18584 15424 18612
rect 13780 18572 13786 18584
rect 15746 18572 15752 18624
rect 15804 18572 15810 18624
rect 1104 18522 18860 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 18860 18522
rect 1104 18448 18860 18470
rect 5626 18408 5632 18420
rect 2746 18380 5632 18408
rect 1394 18164 1400 18216
rect 1452 18164 1458 18216
rect 1673 18207 1731 18213
rect 1673 18173 1685 18207
rect 1719 18204 1731 18207
rect 2746 18204 2774 18380
rect 5626 18368 5632 18380
rect 5684 18368 5690 18420
rect 6454 18368 6460 18420
rect 6512 18368 6518 18420
rect 10226 18368 10232 18420
rect 10284 18408 10290 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 10284 18380 10793 18408
rect 10284 18368 10290 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 10781 18371 10839 18377
rect 12066 18368 12072 18420
rect 12124 18368 12130 18420
rect 13078 18408 13084 18420
rect 12728 18380 13084 18408
rect 4614 18300 4620 18352
rect 4672 18300 4678 18352
rect 6086 18340 6092 18352
rect 5842 18312 6092 18340
rect 6086 18300 6092 18312
rect 6144 18300 6150 18352
rect 11514 18340 11520 18352
rect 10520 18312 11520 18340
rect 4249 18275 4307 18281
rect 4249 18241 4261 18275
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 1719 18176 2774 18204
rect 4264 18204 4292 18235
rect 4338 18232 4344 18284
rect 4396 18232 4402 18284
rect 6178 18232 6184 18284
rect 6236 18272 6242 18284
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 6236 18244 6561 18272
rect 6236 18232 6242 18244
rect 6549 18241 6561 18244
rect 6595 18272 6607 18275
rect 7742 18272 7748 18284
rect 6595 18244 7748 18272
rect 6595 18241 6607 18244
rect 6549 18235 6607 18241
rect 7742 18232 7748 18244
rect 7800 18232 7806 18284
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18272 9459 18275
rect 9858 18272 9864 18284
rect 9447 18244 9864 18272
rect 9447 18241 9459 18244
rect 9401 18235 9459 18241
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 10520 18281 10548 18312
rect 11514 18300 11520 18312
rect 11572 18300 11578 18352
rect 11882 18300 11888 18352
rect 11940 18300 11946 18352
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18241 10563 18275
rect 10505 18235 10563 18241
rect 10686 18232 10692 18284
rect 10744 18232 10750 18284
rect 10965 18275 11023 18281
rect 10965 18241 10977 18275
rect 11011 18272 11023 18275
rect 11146 18272 11152 18284
rect 11011 18244 11152 18272
rect 11011 18241 11023 18244
rect 10965 18235 11023 18241
rect 11146 18232 11152 18244
rect 11204 18232 11210 18284
rect 12728 18281 12756 18380
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 13446 18368 13452 18420
rect 13504 18408 13510 18420
rect 14274 18408 14280 18420
rect 13504 18380 14280 18408
rect 13504 18368 13510 18380
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 14753 18411 14811 18417
rect 14753 18408 14765 18411
rect 14424 18380 14765 18408
rect 14424 18368 14430 18380
rect 14753 18377 14765 18380
rect 14799 18408 14811 18411
rect 15010 18408 15016 18420
rect 14799 18380 15016 18408
rect 14799 18377 14811 18380
rect 14753 18371 14811 18377
rect 15010 18368 15016 18380
rect 15068 18368 15074 18420
rect 12805 18343 12863 18349
rect 12805 18309 12817 18343
rect 12851 18340 12863 18343
rect 12894 18340 12900 18352
rect 12851 18312 12900 18340
rect 12851 18309 12863 18312
rect 12805 18303 12863 18309
rect 12894 18300 12900 18312
rect 12952 18340 12958 18352
rect 13633 18343 13691 18349
rect 13633 18340 13645 18343
rect 12952 18312 13645 18340
rect 12952 18300 12958 18312
rect 13633 18309 13645 18312
rect 13679 18309 13691 18343
rect 13633 18303 13691 18309
rect 14553 18343 14611 18349
rect 14553 18309 14565 18343
rect 14599 18340 14611 18343
rect 15470 18340 15476 18352
rect 14599 18312 15476 18340
rect 14599 18309 14611 18312
rect 14553 18303 14611 18309
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18272 12403 18275
rect 12713 18275 12771 18281
rect 12713 18272 12725 18275
rect 12391 18244 12725 18272
rect 12391 18241 12403 18244
rect 12345 18235 12403 18241
rect 12713 18241 12725 18244
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18241 13047 18275
rect 12989 18235 13047 18241
rect 5350 18204 5356 18216
rect 4264 18176 5356 18204
rect 1719 18173 1731 18176
rect 1673 18167 1731 18173
rect 5350 18164 5356 18176
rect 5408 18164 5414 18216
rect 11241 18207 11299 18213
rect 11241 18173 11253 18207
rect 11287 18204 11299 18207
rect 11698 18204 11704 18216
rect 11287 18176 11704 18204
rect 11287 18173 11299 18176
rect 11241 18167 11299 18173
rect 11698 18164 11704 18176
rect 11756 18204 11762 18216
rect 13004 18204 13032 18235
rect 13446 18232 13452 18284
rect 13504 18232 13510 18284
rect 13722 18232 13728 18284
rect 13780 18232 13786 18284
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14093 18275 14151 18281
rect 14093 18272 14105 18275
rect 13872 18244 14105 18272
rect 13872 18232 13878 18244
rect 14093 18241 14105 18244
rect 14139 18241 14151 18275
rect 14826 18272 14832 18284
rect 14093 18235 14151 18241
rect 14200 18244 14832 18272
rect 14200 18204 14228 18244
rect 14826 18232 14832 18244
rect 14884 18272 14890 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 14884 18244 15209 18272
rect 14884 18232 14890 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 15197 18235 15255 18241
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15381 18275 15439 18281
rect 15381 18272 15393 18275
rect 15344 18244 15393 18272
rect 15344 18232 15350 18244
rect 15381 18241 15393 18244
rect 15427 18241 15439 18275
rect 15381 18235 15439 18241
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 16117 18207 16175 18213
rect 16117 18204 16129 18207
rect 11756 18176 14228 18204
rect 14936 18176 16129 18204
rect 11756 18164 11762 18176
rect 10689 18139 10747 18145
rect 10689 18105 10701 18139
rect 10735 18136 10747 18139
rect 11149 18139 11207 18145
rect 11149 18136 11161 18139
rect 10735 18108 11161 18136
rect 10735 18105 10747 18108
rect 10689 18099 10747 18105
rect 11149 18105 11161 18108
rect 11195 18136 11207 18139
rect 11517 18139 11575 18145
rect 11517 18136 11529 18139
rect 11195 18108 11529 18136
rect 11195 18105 11207 18108
rect 11149 18099 11207 18105
rect 11517 18105 11529 18108
rect 11563 18105 11575 18139
rect 11517 18099 11575 18105
rect 12989 18139 13047 18145
rect 12989 18105 13001 18139
rect 13035 18136 13047 18139
rect 13446 18136 13452 18148
rect 13035 18108 13452 18136
rect 13035 18105 13047 18108
rect 12989 18099 13047 18105
rect 13446 18096 13452 18108
rect 13504 18096 13510 18148
rect 14936 18145 14964 18176
rect 16117 18173 16129 18176
rect 16163 18173 16175 18207
rect 16117 18167 16175 18173
rect 14921 18139 14979 18145
rect 14921 18105 14933 18139
rect 14967 18105 14979 18139
rect 14921 18099 14979 18105
rect 15930 18096 15936 18148
rect 15988 18136 15994 18148
rect 16393 18139 16451 18145
rect 16393 18136 16405 18139
rect 15988 18108 16405 18136
rect 15988 18096 15994 18108
rect 16393 18105 16405 18108
rect 16439 18105 16451 18139
rect 16393 18099 16451 18105
rect 4157 18071 4215 18077
rect 4157 18037 4169 18071
rect 4203 18068 4215 18071
rect 4706 18068 4712 18080
rect 4203 18040 4712 18068
rect 4203 18037 4215 18040
rect 4157 18031 4215 18037
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 5350 18028 5356 18080
rect 5408 18068 5414 18080
rect 6089 18071 6147 18077
rect 6089 18068 6101 18071
rect 5408 18040 6101 18068
rect 5408 18028 5414 18040
rect 6089 18037 6101 18040
rect 6135 18037 6147 18071
rect 6089 18031 6147 18037
rect 9490 18028 9496 18080
rect 9548 18028 9554 18080
rect 11238 18028 11244 18080
rect 11296 18068 11302 18080
rect 11885 18071 11943 18077
rect 11885 18068 11897 18071
rect 11296 18040 11897 18068
rect 11296 18028 11302 18040
rect 11885 18037 11897 18040
rect 11931 18037 11943 18071
rect 11885 18031 11943 18037
rect 12250 18028 12256 18080
rect 12308 18028 12314 18080
rect 13354 18028 13360 18080
rect 13412 18028 13418 18080
rect 13538 18028 13544 18080
rect 13596 18068 13602 18080
rect 14737 18071 14795 18077
rect 14737 18068 14749 18071
rect 13596 18040 14749 18068
rect 13596 18028 13602 18040
rect 14737 18037 14749 18040
rect 14783 18068 14795 18071
rect 15562 18068 15568 18080
rect 14783 18040 15568 18068
rect 14783 18037 14795 18040
rect 14737 18031 14795 18037
rect 15562 18028 15568 18040
rect 15620 18028 15626 18080
rect 1104 17978 18860 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 18860 17978
rect 1104 17904 18860 17926
rect 2590 17824 2596 17876
rect 2648 17824 2654 17876
rect 5169 17867 5227 17873
rect 5169 17833 5181 17867
rect 5215 17864 5227 17867
rect 5258 17864 5264 17876
rect 5215 17836 5264 17864
rect 5215 17833 5227 17836
rect 5169 17827 5227 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 5353 17867 5411 17873
rect 5353 17833 5365 17867
rect 5399 17833 5411 17867
rect 5353 17827 5411 17833
rect 4062 17756 4068 17808
rect 4120 17796 4126 17808
rect 4525 17799 4583 17805
rect 4525 17796 4537 17799
rect 4120 17768 4537 17796
rect 4120 17756 4126 17768
rect 4525 17765 4537 17768
rect 4571 17796 4583 17799
rect 5368 17796 5396 17827
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 6641 17867 6699 17873
rect 6641 17864 6653 17867
rect 6236 17836 6653 17864
rect 6236 17824 6242 17836
rect 6641 17833 6653 17836
rect 6687 17833 6699 17867
rect 6641 17827 6699 17833
rect 10502 17824 10508 17876
rect 10560 17864 10566 17876
rect 11057 17867 11115 17873
rect 11057 17864 11069 17867
rect 10560 17836 11069 17864
rect 10560 17824 10566 17836
rect 11057 17833 11069 17836
rect 11103 17833 11115 17867
rect 11057 17827 11115 17833
rect 11425 17867 11483 17873
rect 11425 17833 11437 17867
rect 11471 17864 11483 17867
rect 11882 17864 11888 17876
rect 11471 17836 11888 17864
rect 11471 17833 11483 17836
rect 11425 17827 11483 17833
rect 11882 17824 11888 17836
rect 11940 17824 11946 17876
rect 4571 17768 5396 17796
rect 4571 17765 4583 17768
rect 4525 17759 4583 17765
rect 14918 17756 14924 17808
rect 14976 17756 14982 17808
rect 15565 17799 15623 17805
rect 15565 17765 15577 17799
rect 15611 17796 15623 17799
rect 15838 17796 15844 17808
rect 15611 17768 15844 17796
rect 15611 17765 15623 17768
rect 15565 17759 15623 17765
rect 15838 17756 15844 17768
rect 15896 17756 15902 17808
rect 2685 17731 2743 17737
rect 2685 17697 2697 17731
rect 2731 17728 2743 17731
rect 2866 17728 2872 17740
rect 2731 17700 2872 17728
rect 2731 17697 2743 17700
rect 2685 17691 2743 17697
rect 2866 17688 2872 17700
rect 2924 17728 2930 17740
rect 3970 17728 3976 17740
rect 2924 17700 3976 17728
rect 2924 17688 2930 17700
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 4448 17700 4936 17728
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2832 17632 2973 17660
rect 2832 17620 2838 17632
rect 2961 17629 2973 17632
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 3142 17620 3148 17672
rect 3200 17620 3206 17672
rect 4448 17669 4476 17700
rect 4908 17669 4936 17700
rect 5350 17688 5356 17740
rect 5408 17688 5414 17740
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 10778 17728 10784 17740
rect 10100 17700 10784 17728
rect 10100 17688 10106 17700
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 15746 17728 15752 17740
rect 15212 17700 15752 17728
rect 4433 17663 4491 17669
rect 4433 17629 4445 17663
rect 4479 17629 4491 17663
rect 4433 17623 4491 17629
rect 4617 17663 4675 17669
rect 4617 17629 4629 17663
rect 4663 17660 4675 17663
rect 4893 17663 4951 17669
rect 4663 17632 4752 17660
rect 4663 17629 4675 17632
rect 4617 17623 4675 17629
rect 4724 17601 4752 17632
rect 4893 17629 4905 17663
rect 4939 17660 4951 17663
rect 5368 17660 5396 17688
rect 4939 17632 5396 17660
rect 4939 17629 4951 17632
rect 4893 17623 4951 17629
rect 6270 17620 6276 17672
rect 6328 17620 6334 17672
rect 11333 17663 11391 17669
rect 11333 17660 11345 17663
rect 11072 17632 11345 17660
rect 4709 17595 4767 17601
rect 4709 17561 4721 17595
rect 4755 17561 4767 17595
rect 4709 17555 4767 17561
rect 5077 17595 5135 17601
rect 5077 17561 5089 17595
rect 5123 17592 5135 17595
rect 5321 17595 5379 17601
rect 5321 17592 5333 17595
rect 5123 17564 5333 17592
rect 5123 17561 5135 17564
rect 5077 17555 5135 17561
rect 5321 17561 5333 17564
rect 5367 17561 5379 17595
rect 5321 17555 5379 17561
rect 5537 17595 5595 17601
rect 5537 17561 5549 17595
rect 5583 17592 5595 17595
rect 5583 17564 6500 17592
rect 5583 17561 5595 17564
rect 5537 17555 5595 17561
rect 2406 17484 2412 17536
rect 2464 17484 2470 17536
rect 2498 17484 2504 17536
rect 2556 17524 2562 17536
rect 2961 17527 3019 17533
rect 2961 17524 2973 17527
rect 2556 17496 2973 17524
rect 2556 17484 2562 17496
rect 2961 17493 2973 17496
rect 3007 17493 3019 17527
rect 4724 17524 4752 17555
rect 6472 17536 6500 17564
rect 9490 17552 9496 17604
rect 9548 17552 9554 17604
rect 10505 17595 10563 17601
rect 10505 17561 10517 17595
rect 10551 17561 10563 17595
rect 10505 17555 10563 17561
rect 5718 17524 5724 17536
rect 4724 17496 5724 17524
rect 2961 17487 3019 17493
rect 5718 17484 5724 17496
rect 5776 17484 5782 17536
rect 6454 17484 6460 17536
rect 6512 17524 6518 17536
rect 6641 17527 6699 17533
rect 6641 17524 6653 17527
rect 6512 17496 6653 17524
rect 6512 17484 6518 17496
rect 6641 17493 6653 17496
rect 6687 17493 6699 17527
rect 6641 17487 6699 17493
rect 6825 17527 6883 17533
rect 6825 17493 6837 17527
rect 6871 17524 6883 17527
rect 7098 17524 7104 17536
rect 6871 17496 7104 17524
rect 6871 17493 6883 17496
rect 6825 17487 6883 17493
rect 7098 17484 7104 17496
rect 7156 17484 7162 17536
rect 9033 17527 9091 17533
rect 9033 17493 9045 17527
rect 9079 17524 9091 17527
rect 10318 17524 10324 17536
rect 9079 17496 10324 17524
rect 9079 17493 9091 17496
rect 9033 17487 9091 17493
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 10520 17524 10548 17555
rect 10594 17552 10600 17604
rect 10652 17592 10658 17604
rect 11072 17601 11100 17632
rect 11333 17629 11345 17632
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 11514 17620 11520 17672
rect 11572 17660 11578 17672
rect 12250 17660 12256 17672
rect 11572 17632 12256 17660
rect 11572 17620 11578 17632
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 14240 17632 14289 17660
rect 14240 17620 14246 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14277 17623 14335 17629
rect 14826 17620 14832 17672
rect 14884 17660 14890 17672
rect 15212 17669 15240 17700
rect 15746 17688 15752 17700
rect 15804 17688 15810 17740
rect 14921 17663 14979 17669
rect 14921 17660 14933 17663
rect 14884 17632 14933 17660
rect 14884 17620 14890 17632
rect 14921 17629 14933 17632
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 15197 17663 15255 17669
rect 15197 17629 15209 17663
rect 15243 17629 15255 17663
rect 15197 17623 15255 17629
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17660 15439 17663
rect 15470 17660 15476 17672
rect 15427 17632 15476 17660
rect 15427 17629 15439 17632
rect 15381 17623 15439 17629
rect 11025 17595 11100 17601
rect 11025 17592 11037 17595
rect 10652 17564 11037 17592
rect 10652 17552 10658 17564
rect 11025 17561 11037 17564
rect 11071 17564 11100 17595
rect 11071 17561 11083 17564
rect 11025 17555 11083 17561
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 11241 17595 11299 17601
rect 11241 17592 11253 17595
rect 11204 17564 11253 17592
rect 11204 17552 11210 17564
rect 11241 17561 11253 17564
rect 11287 17561 11299 17595
rect 11241 17555 11299 17561
rect 15010 17552 15016 17604
rect 15068 17592 15074 17604
rect 15304 17592 15332 17623
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15562 17620 15568 17672
rect 15620 17620 15626 17672
rect 15068 17564 15332 17592
rect 15068 17552 15074 17564
rect 10873 17527 10931 17533
rect 10873 17524 10885 17527
rect 10520 17496 10885 17524
rect 10873 17493 10885 17496
rect 10919 17493 10931 17527
rect 10873 17487 10931 17493
rect 14185 17527 14243 17533
rect 14185 17493 14197 17527
rect 14231 17524 14243 17527
rect 14274 17524 14280 17536
rect 14231 17496 14280 17524
rect 14231 17493 14243 17496
rect 14185 17487 14243 17493
rect 14274 17484 14280 17496
rect 14332 17484 14338 17536
rect 15105 17527 15163 17533
rect 15105 17493 15117 17527
rect 15151 17524 15163 17527
rect 15286 17524 15292 17536
rect 15151 17496 15292 17524
rect 15151 17493 15163 17496
rect 15105 17487 15163 17493
rect 15286 17484 15292 17496
rect 15344 17484 15350 17536
rect 1104 17434 18860 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 18860 17434
rect 1104 17360 18860 17382
rect 2225 17323 2283 17329
rect 2225 17289 2237 17323
rect 2271 17320 2283 17323
rect 2406 17320 2412 17332
rect 2271 17292 2412 17320
rect 2271 17289 2283 17292
rect 2225 17283 2283 17289
rect 2406 17280 2412 17292
rect 2464 17280 2470 17332
rect 3142 17280 3148 17332
rect 3200 17280 3206 17332
rect 4062 17280 4068 17332
rect 4120 17280 4126 17332
rect 5350 17280 5356 17332
rect 5408 17320 5414 17332
rect 5813 17323 5871 17329
rect 5813 17320 5825 17323
rect 5408 17292 5825 17320
rect 5408 17280 5414 17292
rect 5813 17289 5825 17292
rect 5859 17289 5871 17323
rect 5813 17283 5871 17289
rect 6178 17280 6184 17332
rect 6236 17280 6242 17332
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 7800 17292 8984 17320
rect 7800 17280 7806 17292
rect 1673 17255 1731 17261
rect 1673 17221 1685 17255
rect 1719 17252 1731 17255
rect 1762 17252 1768 17264
rect 1719 17224 1768 17252
rect 1719 17221 1731 17224
rect 1673 17215 1731 17221
rect 1762 17212 1768 17224
rect 1820 17212 1826 17264
rect 1889 17255 1947 17261
rect 1889 17221 1901 17255
rect 1935 17252 1947 17255
rect 2498 17252 2504 17264
rect 1935 17224 2504 17252
rect 1935 17221 1947 17224
rect 1889 17215 1947 17221
rect 2148 17193 2176 17224
rect 2498 17212 2504 17224
rect 2556 17212 2562 17264
rect 2593 17255 2651 17261
rect 2593 17221 2605 17255
rect 2639 17252 2651 17255
rect 2961 17255 3019 17261
rect 2961 17252 2973 17255
rect 2639 17224 2973 17252
rect 2639 17221 2651 17224
rect 2593 17215 2651 17221
rect 2961 17221 2973 17224
rect 3007 17221 3019 17255
rect 3160 17252 3188 17280
rect 3160 17224 3740 17252
rect 2961 17215 3019 17221
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2133 17147 2191 17153
rect 2314 17144 2320 17196
rect 2372 17184 2378 17196
rect 2409 17187 2467 17193
rect 2409 17184 2421 17187
rect 2372 17156 2421 17184
rect 2372 17144 2378 17156
rect 2409 17153 2421 17156
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2685 17187 2743 17193
rect 2685 17153 2697 17187
rect 2731 17153 2743 17187
rect 2685 17147 2743 17153
rect 2833 17187 2891 17193
rect 2833 17153 2845 17187
rect 2879 17184 2891 17187
rect 2879 17156 3004 17184
rect 2879 17153 2891 17156
rect 2833 17147 2891 17153
rect 2700 17116 2728 17147
rect 2056 17088 2728 17116
rect 2976 17116 3004 17156
rect 3050 17144 3056 17196
rect 3108 17144 3114 17196
rect 3234 17193 3240 17196
rect 3191 17187 3240 17193
rect 3191 17153 3203 17187
rect 3237 17153 3240 17187
rect 3191 17147 3240 17153
rect 3234 17144 3240 17147
rect 3292 17144 3298 17196
rect 3712 17193 3740 17224
rect 3970 17212 3976 17264
rect 4028 17252 4034 17264
rect 7006 17252 7012 17264
rect 4028 17224 7012 17252
rect 4028 17212 4034 17224
rect 4172 17193 4200 17224
rect 7006 17212 7012 17224
rect 7064 17212 7070 17264
rect 7098 17212 7104 17264
rect 7156 17212 7162 17264
rect 8849 17255 8907 17261
rect 8849 17252 8861 17255
rect 8326 17224 8861 17252
rect 8849 17221 8861 17224
rect 8895 17221 8907 17255
rect 8849 17215 8907 17221
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 3697 17147 3755 17153
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17153 4215 17187
rect 4157 17147 4215 17153
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4798 17184 4804 17196
rect 4479 17156 4804 17184
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 5718 17144 5724 17196
rect 5776 17144 5782 17196
rect 5997 17187 6055 17193
rect 5997 17153 6009 17187
rect 6043 17184 6055 17187
rect 6086 17184 6092 17196
rect 6043 17156 6092 17184
rect 6043 17153 6055 17156
rect 5997 17147 6055 17153
rect 6086 17144 6092 17156
rect 6144 17144 6150 17196
rect 6730 17144 6736 17196
rect 6788 17184 6794 17196
rect 8956 17193 8984 17292
rect 10502 17280 10508 17332
rect 10560 17280 10566 17332
rect 10686 17280 10692 17332
rect 10744 17280 10750 17332
rect 15102 17280 15108 17332
rect 15160 17320 15166 17332
rect 15160 17292 16252 17320
rect 15160 17280 15166 17292
rect 10318 17212 10324 17264
rect 10376 17252 10382 17264
rect 10376 17224 13216 17252
rect 10376 17212 10382 17224
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6788 17156 6837 17184
rect 6788 17144 6794 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9585 17187 9643 17193
rect 9585 17184 9597 17187
rect 9364 17156 9597 17184
rect 9364 17144 9370 17156
rect 9585 17153 9597 17156
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10796 17193 10824 17224
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 10008 17156 10149 17184
rect 10008 17144 10014 17156
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17153 10839 17187
rect 10781 17147 10839 17153
rect 3421 17119 3479 17125
rect 3421 17116 3433 17119
rect 2976 17088 3433 17116
rect 2056 17057 2084 17088
rect 3421 17085 3433 17088
rect 3467 17085 3479 17119
rect 3421 17079 3479 17085
rect 3605 17119 3663 17125
rect 3605 17085 3617 17119
rect 3651 17085 3663 17119
rect 3605 17079 3663 17085
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 4614 17116 4620 17128
rect 4571 17088 4620 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 2041 17051 2099 17057
rect 2041 17017 2053 17051
rect 2087 17017 2099 17051
rect 3620 17048 3648 17079
rect 4614 17076 4620 17088
rect 4672 17076 4678 17128
rect 6104 17116 6132 17144
rect 8573 17119 8631 17125
rect 8573 17116 8585 17119
rect 6104 17088 8585 17116
rect 8573 17085 8585 17088
rect 8619 17085 8631 17119
rect 10152 17116 10180 17147
rect 10612 17116 10640 17147
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 13188 17193 13216 17224
rect 14384 17224 16068 17252
rect 14384 17196 14412 17224
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 10152 17088 10640 17116
rect 12713 17119 12771 17125
rect 8573 17079 8631 17085
rect 12713 17085 12725 17119
rect 12759 17116 12771 17119
rect 12802 17116 12808 17128
rect 12759 17088 12808 17116
rect 12759 17085 12771 17088
rect 12713 17079 12771 17085
rect 12802 17076 12808 17088
rect 12860 17076 12866 17128
rect 13188 17116 13216 17147
rect 13354 17144 13360 17196
rect 13412 17144 13418 17196
rect 14366 17144 14372 17196
rect 14424 17144 14430 17196
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 14507 17156 14596 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 13188 17088 13768 17116
rect 4341 17051 4399 17057
rect 4341 17048 4353 17051
rect 3620 17020 4353 17048
rect 2041 17011 2099 17017
rect 4341 17017 4353 17020
rect 4387 17017 4399 17051
rect 4341 17011 4399 17017
rect 12434 17008 12440 17060
rect 12492 17048 12498 17060
rect 12529 17051 12587 17057
rect 12529 17048 12541 17051
rect 12492 17020 12541 17048
rect 12492 17008 12498 17020
rect 12529 17017 12541 17020
rect 12575 17048 12587 17051
rect 12989 17051 13047 17057
rect 12989 17048 13001 17051
rect 12575 17020 13001 17048
rect 12575 17017 12587 17020
rect 12529 17011 12587 17017
rect 12989 17017 13001 17020
rect 13035 17017 13047 17051
rect 12989 17011 13047 17017
rect 13740 16992 13768 17088
rect 1857 16983 1915 16989
rect 1857 16949 1869 16983
rect 1903 16980 1915 16983
rect 1946 16980 1952 16992
rect 1903 16952 1952 16980
rect 1903 16949 1915 16952
rect 1857 16943 1915 16949
rect 1946 16940 1952 16952
rect 2004 16980 2010 16992
rect 2406 16980 2412 16992
rect 2004 16952 2412 16980
rect 2004 16940 2010 16952
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 3326 16940 3332 16992
rect 3384 16940 3390 16992
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 4706 16980 4712 16992
rect 4295 16952 4712 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 4706 16940 4712 16952
rect 4764 16940 4770 16992
rect 9858 16940 9864 16992
rect 9916 16940 9922 16992
rect 12710 16940 12716 16992
rect 12768 16940 12774 16992
rect 12805 16983 12863 16989
rect 12805 16949 12817 16983
rect 12851 16980 12863 16983
rect 13078 16980 13084 16992
rect 12851 16952 13084 16980
rect 12851 16949 12863 16952
rect 12805 16943 12863 16949
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 14568 16980 14596 17156
rect 14642 17144 14648 17196
rect 14700 17144 14706 17196
rect 14734 17144 14740 17196
rect 14792 17144 14798 17196
rect 14826 17144 14832 17196
rect 14884 17144 14890 17196
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 15120 17193 15148 17224
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 15105 17147 15163 17153
rect 15212 17156 15577 17184
rect 15212 17116 15240 17156
rect 15565 17153 15577 17156
rect 15611 17153 15623 17187
rect 15565 17147 15623 17153
rect 15841 17187 15899 17193
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 15930 17184 15936 17196
rect 15887 17156 15936 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 15930 17144 15936 17156
rect 15988 17144 15994 17196
rect 16040 17193 16068 17224
rect 16224 17193 16252 17292
rect 16025 17187 16083 17193
rect 16025 17153 16037 17187
rect 16071 17153 16083 17187
rect 16025 17147 16083 17153
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 14844 17088 15240 17116
rect 14645 17051 14703 17057
rect 14645 17017 14657 17051
rect 14691 17048 14703 17051
rect 14844 17048 14872 17088
rect 15470 17076 15476 17128
rect 15528 17116 15534 17128
rect 15657 17119 15715 17125
rect 15657 17116 15669 17119
rect 15528 17088 15669 17116
rect 15528 17076 15534 17088
rect 15657 17085 15669 17088
rect 15703 17116 15715 17119
rect 16117 17119 16175 17125
rect 16117 17116 16129 17119
rect 15703 17088 16129 17116
rect 15703 17085 15715 17088
rect 15657 17079 15715 17085
rect 16117 17085 16129 17088
rect 16163 17085 16175 17119
rect 16117 17079 16175 17085
rect 14691 17020 14872 17048
rect 15289 17051 15347 17057
rect 14691 17017 14703 17020
rect 14645 17011 14703 17017
rect 15289 17017 15301 17051
rect 15335 17048 15347 17051
rect 15562 17048 15568 17060
rect 15335 17020 15568 17048
rect 15335 17017 15347 17020
rect 15289 17011 15347 17017
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 15749 17051 15807 17057
rect 15749 17017 15761 17051
rect 15795 17048 15807 17051
rect 15838 17048 15844 17060
rect 15795 17020 15844 17048
rect 15795 17017 15807 17020
rect 15749 17011 15807 17017
rect 15838 17008 15844 17020
rect 15896 17008 15902 17060
rect 15010 16980 15016 16992
rect 13780 16952 15016 16980
rect 13780 16940 13786 16952
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 15378 16940 15384 16992
rect 15436 16940 15442 16992
rect 1104 16890 18860 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 18860 16890
rect 1104 16816 18860 16838
rect 2501 16779 2559 16785
rect 2501 16745 2513 16779
rect 2547 16776 2559 16779
rect 2590 16776 2596 16788
rect 2547 16748 2596 16776
rect 2547 16745 2559 16748
rect 2501 16739 2559 16745
rect 2590 16736 2596 16748
rect 2648 16776 2654 16788
rect 3053 16779 3111 16785
rect 2648 16748 2774 16776
rect 2648 16736 2654 16748
rect 2746 16708 2774 16748
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 3142 16776 3148 16788
rect 3099 16748 3148 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 3142 16736 3148 16748
rect 3200 16736 3206 16788
rect 5445 16779 5503 16785
rect 5445 16776 5457 16779
rect 4908 16748 5457 16776
rect 2746 16680 2912 16708
rect 2409 16643 2467 16649
rect 2409 16609 2421 16643
rect 2455 16640 2467 16643
rect 2884 16640 2912 16680
rect 2455 16612 2774 16640
rect 2884 16612 3004 16640
rect 2455 16609 2467 16612
rect 2409 16603 2467 16609
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16541 1823 16575
rect 1765 16535 1823 16541
rect 1670 16464 1676 16516
rect 1728 16504 1734 16516
rect 1780 16504 1808 16535
rect 1946 16532 1952 16584
rect 2004 16532 2010 16584
rect 2630 16575 2688 16581
rect 2630 16572 2642 16575
rect 2056 16544 2642 16572
rect 2056 16504 2084 16544
rect 2630 16541 2642 16544
rect 2676 16541 2688 16575
rect 2746 16572 2774 16612
rect 2866 16572 2872 16584
rect 2746 16544 2872 16572
rect 2630 16535 2688 16541
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 2976 16572 3004 16612
rect 3421 16575 3479 16581
rect 3421 16572 3433 16575
rect 2976 16544 3433 16572
rect 3421 16541 3433 16544
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 1728 16476 2084 16504
rect 1728 16464 1734 16476
rect 2774 16464 2780 16516
rect 2832 16464 2838 16516
rect 2884 16504 2912 16532
rect 3237 16507 3295 16513
rect 3237 16504 3249 16507
rect 2884 16476 3249 16504
rect 3237 16473 3249 16476
rect 3283 16473 3295 16507
rect 3237 16467 3295 16473
rect 4448 16504 4476 16535
rect 4614 16532 4620 16584
rect 4672 16572 4678 16584
rect 4908 16581 4936 16748
rect 5445 16745 5457 16748
rect 5491 16776 5503 16779
rect 5534 16776 5540 16788
rect 5491 16748 5540 16776
rect 5491 16745 5503 16748
rect 5445 16739 5503 16745
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 5629 16779 5687 16785
rect 5629 16745 5641 16779
rect 5675 16776 5687 16779
rect 6270 16776 6276 16788
rect 5675 16748 6276 16776
rect 5675 16745 5687 16748
rect 5629 16739 5687 16745
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 10410 16736 10416 16788
rect 10468 16736 10474 16788
rect 13722 16736 13728 16788
rect 13780 16736 13786 16788
rect 14366 16736 14372 16788
rect 14424 16776 14430 16788
rect 14553 16779 14611 16785
rect 14553 16776 14565 16779
rect 14424 16748 14565 16776
rect 14424 16736 14430 16748
rect 14553 16745 14565 16748
rect 14599 16745 14611 16779
rect 14553 16739 14611 16745
rect 5350 16668 5356 16720
rect 5408 16708 5414 16720
rect 5721 16711 5779 16717
rect 5721 16708 5733 16711
rect 5408 16680 5733 16708
rect 5408 16668 5414 16680
rect 5721 16677 5733 16680
rect 5767 16677 5779 16711
rect 5721 16671 5779 16677
rect 12253 16711 12311 16717
rect 12253 16677 12265 16711
rect 12299 16708 12311 16711
rect 12437 16711 12495 16717
rect 12437 16708 12449 16711
rect 12299 16680 12449 16708
rect 12299 16677 12311 16680
rect 12253 16671 12311 16677
rect 12437 16677 12449 16680
rect 12483 16677 12495 16711
rect 12437 16671 12495 16677
rect 12728 16680 13952 16708
rect 6638 16640 6644 16652
rect 5184 16612 6644 16640
rect 5184 16581 5212 16612
rect 6638 16600 6644 16612
rect 6696 16600 6702 16652
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12728 16640 12756 16680
rect 11931 16612 12756 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 12802 16600 12808 16652
rect 12860 16640 12866 16652
rect 12897 16643 12955 16649
rect 12897 16640 12909 16643
rect 12860 16612 12909 16640
rect 12860 16600 12866 16612
rect 12897 16609 12909 16612
rect 12943 16640 12955 16643
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 12943 16612 13277 16640
rect 12943 16609 12955 16612
rect 12897 16603 12955 16609
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 13354 16600 13360 16652
rect 13412 16640 13418 16652
rect 13412 16612 13676 16640
rect 13412 16600 13418 16612
rect 4801 16575 4859 16581
rect 4801 16572 4813 16575
rect 4672 16544 4813 16572
rect 4672 16532 4678 16544
rect 4801 16541 4813 16544
rect 4847 16541 4859 16575
rect 4801 16535 4859 16541
rect 4893 16575 4951 16581
rect 4893 16541 4905 16575
rect 4939 16541 4951 16575
rect 4893 16535 4951 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 5184 16504 5212 16535
rect 5350 16532 5356 16584
rect 5408 16532 5414 16584
rect 5718 16532 5724 16584
rect 5776 16572 5782 16584
rect 5905 16575 5963 16581
rect 5905 16572 5917 16575
rect 5776 16544 5917 16572
rect 5776 16532 5782 16544
rect 5905 16541 5917 16544
rect 5951 16541 5963 16575
rect 5905 16535 5963 16541
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 6052 16544 6224 16572
rect 6052 16532 6058 16544
rect 4448 16476 5212 16504
rect 5261 16507 5319 16513
rect 1854 16396 1860 16448
rect 1912 16396 1918 16448
rect 2133 16439 2191 16445
rect 2133 16405 2145 16439
rect 2179 16436 2191 16439
rect 2590 16436 2596 16448
rect 2179 16408 2596 16436
rect 2179 16405 2191 16408
rect 2133 16399 2191 16405
rect 2590 16396 2596 16408
rect 2648 16396 2654 16448
rect 2792 16436 2820 16464
rect 4448 16436 4476 16476
rect 5261 16473 5273 16507
rect 5307 16504 5319 16507
rect 5368 16504 5396 16532
rect 5307 16476 5396 16504
rect 5477 16507 5535 16513
rect 5307 16473 5319 16476
rect 5261 16467 5319 16473
rect 5477 16473 5489 16507
rect 5523 16504 5535 16507
rect 6196 16504 6224 16544
rect 6270 16532 6276 16584
rect 6328 16572 6334 16584
rect 6365 16575 6423 16581
rect 6365 16572 6377 16575
rect 6328 16544 6377 16572
rect 6328 16532 6334 16544
rect 6365 16541 6377 16544
rect 6411 16541 6423 16575
rect 11974 16572 11980 16584
rect 6365 16535 6423 16541
rect 10612 16544 11980 16572
rect 6549 16507 6607 16513
rect 6549 16504 6561 16507
rect 5523 16476 6132 16504
rect 6196 16476 6561 16504
rect 5523 16473 5535 16476
rect 5477 16467 5535 16473
rect 6104 16448 6132 16476
rect 6549 16473 6561 16476
rect 6595 16473 6607 16507
rect 6549 16467 6607 16473
rect 9122 16464 9128 16516
rect 9180 16504 9186 16516
rect 10612 16513 10640 16544
rect 11974 16532 11980 16544
rect 12032 16572 12038 16584
rect 12069 16575 12127 16581
rect 12069 16572 12081 16575
rect 12032 16544 12081 16572
rect 12032 16532 12038 16544
rect 12069 16541 12081 16544
rect 12115 16572 12127 16575
rect 13449 16575 13507 16581
rect 13449 16572 13461 16575
rect 12115 16544 13461 16572
rect 12115 16541 12127 16544
rect 12069 16535 12127 16541
rect 13449 16541 13461 16544
rect 13495 16541 13507 16575
rect 13449 16535 13507 16541
rect 13541 16575 13599 16581
rect 13541 16541 13553 16575
rect 13587 16541 13599 16575
rect 13648 16572 13676 16612
rect 13817 16575 13875 16581
rect 13817 16572 13829 16575
rect 13648 16544 13829 16572
rect 13541 16535 13599 16541
rect 13817 16541 13829 16544
rect 13863 16541 13875 16575
rect 13817 16535 13875 16541
rect 10597 16507 10655 16513
rect 9180 16476 10364 16504
rect 9180 16464 9186 16476
rect 2792 16408 4476 16436
rect 4614 16396 4620 16448
rect 4672 16396 4678 16448
rect 5077 16439 5135 16445
rect 5077 16405 5089 16439
rect 5123 16436 5135 16439
rect 5350 16436 5356 16448
rect 5123 16408 5356 16436
rect 5123 16405 5135 16408
rect 5077 16399 5135 16405
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 5994 16396 6000 16448
rect 6052 16396 6058 16448
rect 6086 16396 6092 16448
rect 6144 16396 6150 16448
rect 6270 16396 6276 16448
rect 6328 16396 6334 16448
rect 6638 16396 6644 16448
rect 6696 16436 6702 16448
rect 6733 16439 6791 16445
rect 6733 16436 6745 16439
rect 6696 16408 6745 16436
rect 6696 16396 6702 16408
rect 6733 16405 6745 16408
rect 6779 16405 6791 16439
rect 6733 16399 6791 16405
rect 9950 16396 9956 16448
rect 10008 16436 10014 16448
rect 10229 16439 10287 16445
rect 10229 16436 10241 16439
rect 10008 16408 10241 16436
rect 10008 16396 10014 16408
rect 10229 16405 10241 16408
rect 10275 16405 10287 16439
rect 10336 16436 10364 16476
rect 10597 16473 10609 16507
rect 10643 16473 10655 16507
rect 10597 16467 10655 16473
rect 12434 16464 12440 16516
rect 12492 16464 12498 16516
rect 10397 16439 10455 16445
rect 10397 16436 10409 16439
rect 10336 16408 10409 16436
rect 10229 16399 10287 16405
rect 10397 16405 10409 16408
rect 10443 16436 10455 16439
rect 10870 16436 10876 16448
rect 10443 16408 10876 16436
rect 10443 16405 10455 16408
rect 10397 16399 10455 16405
rect 10870 16396 10876 16408
rect 10928 16396 10934 16448
rect 12986 16396 12992 16448
rect 13044 16396 13050 16448
rect 13170 16396 13176 16448
rect 13228 16396 13234 16448
rect 13464 16436 13492 16535
rect 13556 16504 13584 16535
rect 13924 16504 13952 16680
rect 14369 16643 14427 16649
rect 14369 16609 14381 16643
rect 14415 16640 14427 16643
rect 14550 16640 14556 16652
rect 14415 16612 14556 16640
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 14550 16600 14556 16612
rect 14608 16600 14614 16652
rect 14274 16532 14280 16584
rect 14332 16532 14338 16584
rect 14918 16532 14924 16584
rect 14976 16532 14982 16584
rect 15470 16532 15476 16584
rect 15528 16532 15534 16584
rect 15562 16532 15568 16584
rect 15620 16572 15626 16584
rect 15749 16575 15807 16581
rect 15749 16572 15761 16575
rect 15620 16544 15761 16572
rect 15620 16532 15626 16544
rect 15749 16541 15761 16544
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 15838 16532 15844 16584
rect 15896 16572 15902 16584
rect 16117 16575 16175 16581
rect 16117 16572 16129 16575
rect 15896 16544 16129 16572
rect 15896 16532 15902 16544
rect 16117 16541 16129 16544
rect 16163 16541 16175 16575
rect 16117 16535 16175 16541
rect 14292 16504 14320 16532
rect 13556 16476 14320 16504
rect 14366 16436 14372 16448
rect 13464 16408 14372 16436
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 16117 16439 16175 16445
rect 16117 16405 16129 16439
rect 16163 16436 16175 16439
rect 16206 16436 16212 16448
rect 16163 16408 16212 16436
rect 16163 16405 16175 16408
rect 16117 16399 16175 16405
rect 16206 16396 16212 16408
rect 16264 16396 16270 16448
rect 1104 16346 18860 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 18860 16346
rect 1104 16272 18860 16294
rect 1762 16192 1768 16244
rect 1820 16232 1826 16244
rect 2314 16232 2320 16244
rect 1820 16204 2320 16232
rect 1820 16192 1826 16204
rect 2314 16192 2320 16204
rect 2372 16232 2378 16244
rect 6086 16232 6092 16244
rect 2372 16204 6092 16232
rect 2372 16192 2378 16204
rect 6086 16192 6092 16204
rect 6144 16192 6150 16244
rect 8113 16235 8171 16241
rect 8113 16201 8125 16235
rect 8159 16232 8171 16235
rect 12713 16235 12771 16241
rect 8159 16204 10456 16232
rect 8159 16201 8171 16204
rect 8113 16195 8171 16201
rect 10428 16176 10456 16204
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 12986 16232 12992 16244
rect 12759 16204 12992 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 13262 16192 13268 16244
rect 13320 16192 13326 16244
rect 14384 16204 14688 16232
rect 2041 16167 2099 16173
rect 2041 16133 2053 16167
rect 2087 16164 2099 16167
rect 2682 16164 2688 16176
rect 2087 16136 2688 16164
rect 2087 16133 2099 16136
rect 2041 16127 2099 16133
rect 2682 16124 2688 16136
rect 2740 16164 2746 16176
rect 4798 16164 4804 16176
rect 2740 16136 4804 16164
rect 2740 16124 2746 16136
rect 842 16056 848 16108
rect 900 16096 906 16108
rect 1489 16099 1547 16105
rect 1489 16096 1501 16099
rect 900 16068 1501 16096
rect 900 16056 906 16068
rect 1489 16065 1501 16068
rect 1535 16065 1547 16099
rect 1489 16059 1547 16065
rect 1854 16056 1860 16108
rect 1912 16096 1918 16108
rect 4724 16105 4752 16136
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 4985 16167 5043 16173
rect 4985 16133 4997 16167
rect 5031 16164 5043 16167
rect 5350 16164 5356 16176
rect 5031 16136 5356 16164
rect 5031 16133 5043 16136
rect 4985 16127 5043 16133
rect 5350 16124 5356 16136
rect 5408 16124 5414 16176
rect 6454 16124 6460 16176
rect 6512 16164 6518 16176
rect 6733 16167 6791 16173
rect 6733 16164 6745 16167
rect 6512 16136 6745 16164
rect 6512 16124 6518 16136
rect 6733 16133 6745 16136
rect 6779 16133 6791 16167
rect 6733 16127 6791 16133
rect 9030 16124 9036 16176
rect 9088 16124 9094 16176
rect 10321 16167 10379 16173
rect 10321 16133 10333 16167
rect 10367 16133 10379 16167
rect 10321 16127 10379 16133
rect 2777 16099 2835 16105
rect 2777 16096 2789 16099
rect 1912 16068 2789 16096
rect 1912 16056 1918 16068
rect 2777 16065 2789 16068
rect 2823 16065 2835 16099
rect 2777 16059 2835 16065
rect 4709 16099 4767 16105
rect 4709 16065 4721 16099
rect 4755 16065 4767 16099
rect 4709 16059 4767 16065
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16096 5135 16099
rect 5718 16096 5724 16108
rect 5123 16068 5724 16096
rect 5123 16065 5135 16068
rect 5077 16059 5135 16065
rect 5718 16056 5724 16068
rect 5776 16056 5782 16108
rect 6270 16056 6276 16108
rect 6328 16096 6334 16108
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 6328 16068 6377 16096
rect 6328 16056 6334 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 7742 16056 7748 16108
rect 7800 16056 7806 16108
rect 9861 16099 9919 16105
rect 9861 16065 9873 16099
rect 9907 16096 9919 16099
rect 10042 16096 10048 16108
rect 9907 16068 10048 16096
rect 9907 16065 9919 16068
rect 9861 16059 9919 16065
rect 10042 16056 10048 16068
rect 10100 16056 10106 16108
rect 2590 15988 2596 16040
rect 2648 15988 2654 16040
rect 4617 16031 4675 16037
rect 4617 15997 4629 16031
rect 4663 16028 4675 16031
rect 4890 16028 4896 16040
rect 4663 16000 4896 16028
rect 4663 15997 4675 16000
rect 4617 15991 4675 15997
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 9490 15988 9496 16040
rect 9548 16028 9554 16040
rect 9585 16031 9643 16037
rect 9585 16028 9597 16031
rect 9548 16000 9597 16028
rect 9548 15988 9554 16000
rect 9585 15997 9597 16000
rect 9631 15997 9643 16031
rect 9585 15991 9643 15997
rect 9950 15988 9956 16040
rect 10008 15988 10014 16040
rect 10336 16028 10364 16127
rect 10410 16124 10416 16176
rect 10468 16164 10474 16176
rect 10965 16167 11023 16173
rect 10965 16164 10977 16167
rect 10468 16136 10977 16164
rect 10468 16124 10474 16136
rect 10965 16133 10977 16136
rect 11011 16164 11023 16167
rect 13280 16164 13308 16192
rect 14384 16176 14412 16204
rect 11011 16136 12434 16164
rect 11011 16133 11023 16136
rect 10965 16127 11023 16133
rect 10781 16099 10839 16105
rect 10781 16065 10793 16099
rect 10827 16065 10839 16099
rect 10781 16059 10839 16065
rect 10796 16028 10824 16059
rect 10870 16056 10876 16108
rect 10928 16096 10934 16108
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 10928 16068 11069 16096
rect 10928 16056 10934 16068
rect 11057 16065 11069 16068
rect 11103 16096 11115 16099
rect 11238 16096 11244 16108
rect 11103 16068 11244 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11514 16056 11520 16108
rect 11572 16096 11578 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11572 16068 11713 16096
rect 11572 16056 11578 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11974 16028 11980 16040
rect 10336 16000 10732 16028
rect 10796 16000 11980 16028
rect 3878 15920 3884 15972
rect 3936 15960 3942 15972
rect 5994 15960 6000 15972
rect 3936 15932 6000 15960
rect 3936 15920 3942 15932
rect 5994 15920 6000 15932
rect 6052 15920 6058 15972
rect 10597 15963 10655 15969
rect 10597 15960 10609 15963
rect 10336 15932 10609 15960
rect 2961 15895 3019 15901
rect 2961 15861 2973 15895
rect 3007 15892 3019 15895
rect 3234 15892 3240 15904
rect 3007 15864 3240 15892
rect 3007 15861 3019 15864
rect 2961 15855 3019 15861
rect 3234 15852 3240 15864
rect 3292 15892 3298 15904
rect 3694 15892 3700 15904
rect 3292 15864 3700 15892
rect 3292 15852 3298 15864
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 4433 15895 4491 15901
rect 4433 15861 4445 15895
rect 4479 15892 4491 15895
rect 4798 15892 4804 15904
rect 4479 15864 4804 15892
rect 4479 15861 4491 15864
rect 4433 15855 4491 15861
rect 4798 15852 4804 15864
rect 4856 15852 4862 15904
rect 6638 15852 6644 15904
rect 6696 15892 6702 15904
rect 6733 15895 6791 15901
rect 6733 15892 6745 15895
rect 6696 15864 6745 15892
rect 6696 15852 6702 15864
rect 6733 15861 6745 15864
rect 6779 15861 6791 15895
rect 6733 15855 6791 15861
rect 6914 15852 6920 15904
rect 6972 15852 6978 15904
rect 7650 15852 7656 15904
rect 7708 15852 7714 15904
rect 10336 15901 10364 15932
rect 10597 15929 10609 15932
rect 10643 15929 10655 15963
rect 10704 15960 10732 16000
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 11146 15960 11152 15972
rect 10704 15932 11152 15960
rect 10597 15923 10655 15929
rect 11146 15920 11152 15932
rect 11204 15960 11210 15972
rect 11882 15960 11888 15972
rect 11204 15932 11888 15960
rect 11204 15920 11210 15932
rect 11882 15920 11888 15932
rect 11940 15920 11946 15972
rect 12406 15960 12434 16136
rect 13188 16136 13308 16164
rect 12894 16056 12900 16108
rect 12952 16056 12958 16108
rect 13078 16056 13084 16108
rect 13136 16056 13142 16108
rect 13188 16105 13216 16136
rect 14366 16124 14372 16176
rect 14424 16124 14430 16176
rect 14569 16167 14627 16173
rect 14569 16164 14581 16167
rect 14568 16133 14581 16164
rect 14615 16133 14627 16167
rect 14660 16164 14688 16204
rect 14734 16192 14740 16244
rect 14792 16192 14798 16244
rect 15749 16235 15807 16241
rect 15749 16201 15761 16235
rect 15795 16232 15807 16235
rect 16666 16232 16672 16244
rect 15795 16204 16672 16232
rect 15795 16201 15807 16204
rect 15749 16195 15807 16201
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 15105 16167 15163 16173
rect 15105 16164 15117 16167
rect 14660 16136 15117 16164
rect 14568 16127 14627 16133
rect 15105 16133 15117 16136
rect 15151 16133 15163 16167
rect 15105 16127 15163 16133
rect 13173 16099 13231 16105
rect 13173 16065 13185 16099
rect 13219 16065 13231 16099
rect 13173 16059 13231 16065
rect 13262 16056 13268 16108
rect 13320 16056 13326 16108
rect 13446 16056 13452 16108
rect 13504 16056 13510 16108
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14568 16096 14596 16127
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 15930 16164 15936 16176
rect 15344 16136 15936 16164
rect 15344 16124 15350 16136
rect 15930 16124 15936 16136
rect 15988 16164 15994 16176
rect 15988 16136 16344 16164
rect 15988 16124 15994 16136
rect 14829 16099 14887 16105
rect 14829 16096 14841 16099
rect 14516 16068 14841 16096
rect 14516 16056 14522 16068
rect 14829 16065 14841 16068
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 14918 16056 14924 16108
rect 14976 16056 14982 16108
rect 15378 16056 15384 16108
rect 15436 16056 15442 16108
rect 15808 16099 15866 16105
rect 15808 16065 15820 16099
rect 15854 16096 15866 16099
rect 16025 16099 16083 16105
rect 16025 16096 16037 16099
rect 15854 16068 16037 16096
rect 15854 16065 15866 16068
rect 15808 16059 15866 16065
rect 16025 16065 16037 16068
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 16206 16056 16212 16108
rect 16264 16056 16270 16108
rect 16316 16105 16344 16136
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 15010 15988 15016 16040
rect 15068 16028 15074 16040
rect 15289 16031 15347 16037
rect 15289 16028 15301 16031
rect 15068 16000 15301 16028
rect 15068 15988 15074 16000
rect 15289 15997 15301 16000
rect 15335 15997 15347 16031
rect 15289 15991 15347 15997
rect 13538 15960 13544 15972
rect 12406 15932 13544 15960
rect 13538 15920 13544 15932
rect 13596 15920 13602 15972
rect 15105 15963 15163 15969
rect 15105 15929 15117 15963
rect 15151 15960 15163 15963
rect 15194 15960 15200 15972
rect 15151 15932 15200 15960
rect 15151 15929 15163 15932
rect 15105 15923 15163 15929
rect 15194 15920 15200 15932
rect 15252 15920 15258 15972
rect 10321 15895 10379 15901
rect 10321 15861 10333 15895
rect 10367 15861 10379 15895
rect 10321 15855 10379 15861
rect 10502 15852 10508 15904
rect 10560 15852 10566 15904
rect 11606 15852 11612 15904
rect 11664 15852 11670 15904
rect 14550 15852 14556 15904
rect 14608 15892 14614 15904
rect 14918 15892 14924 15904
rect 14608 15864 14924 15892
rect 14608 15852 14614 15864
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15930 15852 15936 15904
rect 15988 15852 15994 15904
rect 1104 15802 18860 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 18860 15802
rect 1104 15728 18860 15750
rect 4338 15648 4344 15700
rect 4396 15688 4402 15700
rect 4396 15660 5028 15688
rect 4396 15648 4402 15660
rect 4154 15580 4160 15632
rect 4212 15620 4218 15632
rect 4433 15623 4491 15629
rect 4433 15620 4445 15623
rect 4212 15592 4445 15620
rect 4212 15580 4218 15592
rect 4433 15589 4445 15592
rect 4479 15589 4491 15623
rect 4890 15620 4896 15632
rect 4433 15583 4491 15589
rect 4540 15592 4896 15620
rect 1762 15512 1768 15564
rect 1820 15512 1826 15564
rect 2041 15555 2099 15561
rect 2041 15521 2053 15555
rect 2087 15552 2099 15555
rect 2866 15552 2872 15564
rect 2087 15524 2872 15552
rect 2087 15521 2099 15524
rect 2041 15515 2099 15521
rect 2866 15512 2872 15524
rect 2924 15512 2930 15564
rect 4540 15552 4568 15592
rect 4890 15580 4896 15592
rect 4948 15580 4954 15632
rect 4172 15524 4568 15552
rect 1670 15444 1676 15496
rect 1728 15444 1734 15496
rect 2682 15444 2688 15496
rect 2740 15484 2746 15496
rect 4172 15493 4200 15524
rect 4614 15512 4620 15564
rect 4672 15552 4678 15564
rect 4672 15524 4936 15552
rect 4672 15512 4678 15524
rect 3973 15487 4031 15493
rect 3973 15484 3985 15487
rect 2740 15456 3985 15484
rect 2740 15444 2746 15456
rect 3973 15453 3985 15456
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15453 4215 15487
rect 4157 15447 4215 15453
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 4264 15348 4292 15447
rect 4338 15444 4344 15496
rect 4396 15444 4402 15496
rect 4706 15444 4712 15496
rect 4764 15444 4770 15496
rect 4798 15444 4804 15496
rect 4856 15444 4862 15496
rect 4908 15493 4936 15524
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15453 4951 15487
rect 5000 15484 5028 15660
rect 5994 15648 6000 15700
rect 6052 15688 6058 15700
rect 6457 15691 6515 15697
rect 6457 15688 6469 15691
rect 6052 15660 6469 15688
rect 6052 15648 6058 15660
rect 6457 15657 6469 15660
rect 6503 15657 6515 15691
rect 6457 15651 6515 15657
rect 9490 15648 9496 15700
rect 9548 15648 9554 15700
rect 9677 15691 9735 15697
rect 9677 15657 9689 15691
rect 9723 15657 9735 15691
rect 9677 15651 9735 15657
rect 9401 15623 9459 15629
rect 9401 15589 9413 15623
rect 9447 15620 9459 15623
rect 9692 15620 9720 15651
rect 11974 15648 11980 15700
rect 12032 15648 12038 15700
rect 16393 15691 16451 15697
rect 16393 15657 16405 15691
rect 16439 15688 16451 15691
rect 17770 15688 17776 15700
rect 16439 15660 17776 15688
rect 16439 15657 16451 15660
rect 16393 15651 16451 15657
rect 17770 15648 17776 15660
rect 17828 15688 17834 15700
rect 17865 15691 17923 15697
rect 17865 15688 17877 15691
rect 17828 15660 17877 15688
rect 17828 15648 17834 15660
rect 17865 15657 17877 15660
rect 17911 15657 17923 15691
rect 17865 15651 17923 15657
rect 9447 15592 9720 15620
rect 9447 15589 9459 15592
rect 9401 15583 9459 15589
rect 11514 15580 11520 15632
rect 11572 15620 11578 15632
rect 12434 15620 12440 15632
rect 11572 15592 12440 15620
rect 11572 15580 11578 15592
rect 12434 15580 12440 15592
rect 12492 15580 12498 15632
rect 12710 15580 12716 15632
rect 12768 15580 12774 15632
rect 16206 15620 16212 15632
rect 14936 15592 16212 15620
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 6972 15524 7941 15552
rect 6972 15512 6978 15524
rect 7929 15521 7941 15524
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 8205 15555 8263 15561
rect 8205 15521 8217 15555
rect 8251 15552 8263 15555
rect 10042 15552 10048 15564
rect 8251 15524 10048 15552
rect 8251 15521 8263 15524
rect 8205 15515 8263 15521
rect 10042 15512 10048 15524
rect 10100 15552 10106 15564
rect 10229 15555 10287 15561
rect 10229 15552 10241 15555
rect 10100 15524 10241 15552
rect 10100 15512 10106 15524
rect 10229 15521 10241 15524
rect 10275 15521 10287 15555
rect 10229 15515 10287 15521
rect 10502 15512 10508 15564
rect 10560 15512 10566 15564
rect 12728 15552 12756 15580
rect 12728 15524 12940 15552
rect 5077 15487 5135 15493
rect 5077 15484 5089 15487
rect 5000 15456 5089 15484
rect 4893 15447 4951 15453
rect 5077 15453 5089 15456
rect 5123 15453 5135 15487
rect 5077 15447 5135 15453
rect 6089 15487 6147 15493
rect 6089 15453 6101 15487
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 4522 15376 4528 15428
rect 4580 15416 4586 15428
rect 5261 15419 5319 15425
rect 5261 15416 5273 15419
rect 4580 15388 5273 15416
rect 4580 15376 4586 15388
rect 5261 15385 5273 15388
rect 5307 15385 5319 15419
rect 6104 15416 6132 15447
rect 6270 15444 6276 15496
rect 6328 15444 6334 15496
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 9217 15487 9275 15493
rect 9217 15484 9229 15487
rect 8803 15456 9229 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 9217 15453 9229 15456
rect 9263 15484 9275 15487
rect 9263 15456 9996 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 6362 15416 6368 15428
rect 6104 15388 6368 15416
rect 5261 15379 5319 15385
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 7650 15416 7656 15428
rect 7498 15388 7656 15416
rect 7650 15376 7656 15388
rect 7708 15376 7714 15428
rect 8588 15416 8616 15447
rect 9033 15419 9091 15425
rect 9033 15416 9045 15419
rect 8588 15388 9045 15416
rect 9033 15385 9045 15388
rect 9079 15416 9091 15419
rect 9122 15416 9128 15428
rect 9079 15388 9128 15416
rect 9079 15385 9091 15388
rect 9033 15379 9091 15385
rect 9122 15376 9128 15388
rect 9180 15376 9186 15428
rect 9766 15376 9772 15428
rect 9824 15416 9830 15428
rect 9861 15419 9919 15425
rect 9861 15416 9873 15419
rect 9824 15388 9873 15416
rect 9824 15376 9830 15388
rect 9861 15385 9873 15388
rect 9907 15385 9919 15419
rect 9968 15416 9996 15456
rect 11606 15444 11612 15496
rect 11664 15444 11670 15496
rect 12710 15444 12716 15496
rect 12768 15444 12774 15496
rect 12912 15493 12940 15524
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 13081 15487 13139 15493
rect 13081 15453 13093 15487
rect 13127 15484 13139 15487
rect 13446 15484 13452 15496
rect 13127 15456 13452 15484
rect 13127 15453 13139 15456
rect 13081 15447 13139 15453
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 14936 15493 14964 15592
rect 16206 15580 16212 15592
rect 16264 15580 16270 15632
rect 17681 15623 17739 15629
rect 17681 15589 17693 15623
rect 17727 15589 17739 15623
rect 17681 15583 17739 15589
rect 15470 15512 15476 15564
rect 15528 15512 15534 15564
rect 17696 15552 17724 15583
rect 15580 15524 17724 15552
rect 14921 15487 14979 15493
rect 14921 15453 14933 15487
rect 14967 15453 14979 15487
rect 14921 15447 14979 15453
rect 15286 15444 15292 15496
rect 15344 15444 15350 15496
rect 15580 15493 15608 15524
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15453 15623 15487
rect 15565 15447 15623 15453
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15453 16359 15487
rect 16301 15447 16359 15453
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15484 16543 15487
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 16531 15456 17233 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 17221 15453 17233 15456
rect 17267 15484 17279 15487
rect 17310 15484 17316 15496
rect 17267 15456 17316 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 10410 15416 10416 15428
rect 9968 15388 10416 15416
rect 9861 15379 9919 15385
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 12805 15419 12863 15425
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 13170 15416 13176 15428
rect 12851 15388 13176 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 13170 15376 13176 15388
rect 13228 15376 13234 15428
rect 16316 15416 16344 15447
rect 17310 15444 17316 15456
rect 17368 15444 17374 15496
rect 16574 15416 16580 15428
rect 16316 15388 16580 15416
rect 16574 15376 16580 15388
rect 16632 15416 16638 15428
rect 17405 15419 17463 15425
rect 17405 15416 17417 15419
rect 16632 15388 17417 15416
rect 16632 15376 16638 15388
rect 17405 15385 17417 15388
rect 17451 15385 17463 15419
rect 17833 15419 17891 15425
rect 17833 15416 17845 15419
rect 17405 15379 17463 15385
rect 17604 15388 17845 15416
rect 17604 15360 17632 15388
rect 17833 15385 17845 15388
rect 17879 15385 17891 15419
rect 17833 15379 17891 15385
rect 17954 15376 17960 15428
rect 18012 15416 18018 15428
rect 18049 15419 18107 15425
rect 18049 15416 18061 15419
rect 18012 15388 18061 15416
rect 18012 15376 18018 15388
rect 18049 15385 18061 15388
rect 18095 15385 18107 15419
rect 18049 15379 18107 15385
rect 5350 15348 5356 15360
rect 4264 15320 5356 15348
rect 5350 15308 5356 15320
rect 5408 15308 5414 15360
rect 6086 15308 6092 15360
rect 6144 15308 6150 15360
rect 8757 15351 8815 15357
rect 8757 15317 8769 15351
rect 8803 15348 8815 15351
rect 9651 15351 9709 15357
rect 9651 15348 9663 15351
rect 8803 15320 9663 15348
rect 8803 15317 8815 15320
rect 8757 15311 8815 15317
rect 9651 15317 9663 15320
rect 9697 15317 9709 15351
rect 9651 15311 9709 15317
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 12894 15348 12900 15360
rect 12575 15320 12900 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 17586 15308 17592 15360
rect 17644 15308 17650 15360
rect 1104 15258 18860 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 18860 15258
rect 1104 15184 18860 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 1670 15144 1676 15156
rect 1627 15116 1676 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 1670 15104 1676 15116
rect 1728 15104 1734 15156
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15113 2835 15147
rect 2777 15107 2835 15113
rect 3237 15147 3295 15153
rect 3237 15113 3249 15147
rect 3283 15144 3295 15147
rect 4338 15144 4344 15156
rect 3283 15116 4344 15144
rect 3283 15113 3295 15116
rect 3237 15107 3295 15113
rect 842 14968 848 15020
rect 900 15008 906 15020
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 900 14980 1409 15008
rect 900 14968 906 14980
rect 1397 14977 1409 14980
rect 1443 14977 1455 15011
rect 1688 15008 1716 15104
rect 2792 15076 2820 15107
rect 4338 15104 4344 15116
rect 4396 15104 4402 15156
rect 5353 15147 5411 15153
rect 5353 15113 5365 15147
rect 5399 15144 5411 15147
rect 8570 15144 8576 15156
rect 5399 15116 8576 15144
rect 5399 15113 5411 15116
rect 5353 15107 5411 15113
rect 8570 15104 8576 15116
rect 8628 15104 8634 15156
rect 9030 15104 9036 15156
rect 9088 15104 9094 15156
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10870 15144 10876 15156
rect 10100 15116 10876 15144
rect 10100 15104 10106 15116
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 11238 15144 11244 15156
rect 11020 15116 11244 15144
rect 11020 15104 11026 15116
rect 11238 15104 11244 15116
rect 11296 15144 11302 15156
rect 11296 15116 12756 15144
rect 11296 15104 11302 15116
rect 2792 15048 4476 15076
rect 2225 15011 2283 15017
rect 2225 15008 2237 15011
rect 1688 14980 2237 15008
rect 1397 14971 1455 14977
rect 2225 14977 2237 14980
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2866 14968 2872 15020
rect 2924 14968 2930 15020
rect 3326 14968 3332 15020
rect 3384 14968 3390 15020
rect 3510 14968 3516 15020
rect 3568 14968 3574 15020
rect 3694 14968 3700 15020
rect 3752 14968 3758 15020
rect 3878 14968 3884 15020
rect 3936 14968 3942 15020
rect 4448 15017 4476 15048
rect 4614 15036 4620 15088
rect 4672 15036 4678 15088
rect 5810 15036 5816 15088
rect 5868 15036 5874 15088
rect 5994 15036 6000 15088
rect 6052 15085 6058 15088
rect 6052 15079 6071 15085
rect 6059 15045 6071 15079
rect 6730 15076 6736 15088
rect 6052 15039 6071 15045
rect 6380 15048 6736 15076
rect 6052 15036 6058 15039
rect 4433 15011 4491 15017
rect 4433 14977 4445 15011
rect 4479 14977 4491 15011
rect 4433 14971 4491 14977
rect 4522 14968 4528 15020
rect 4580 14968 4586 15020
rect 4632 15008 4660 15036
rect 6380 15017 6408 15048
rect 6730 15036 6736 15048
rect 6788 15036 6794 15088
rect 7650 15036 7656 15088
rect 7708 15036 7714 15088
rect 8757 15079 8815 15085
rect 8757 15045 8769 15079
rect 8803 15076 8815 15079
rect 11330 15076 11336 15088
rect 8803 15048 11336 15076
rect 8803 15045 8815 15048
rect 8757 15039 8815 15045
rect 11330 15036 11336 15048
rect 11388 15076 11394 15088
rect 11388 15048 11744 15076
rect 11388 15036 11394 15048
rect 4801 15011 4859 15017
rect 4801 15008 4813 15011
rect 4632 14980 4813 15008
rect 4801 14977 4813 14980
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 9125 15011 9183 15017
rect 9125 14977 9137 15011
rect 9171 14977 9183 15011
rect 9125 14971 9183 14977
rect 1670 14900 1676 14952
rect 1728 14900 1734 14952
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 2501 14943 2559 14949
rect 2501 14940 2513 14943
rect 1820 14912 2513 14940
rect 1820 14900 1826 14912
rect 2501 14909 2513 14912
rect 2547 14909 2559 14943
rect 2961 14943 3019 14949
rect 2961 14940 2973 14943
rect 2501 14903 2559 14909
rect 2746 14912 2973 14940
rect 2041 14875 2099 14881
rect 2041 14841 2053 14875
rect 2087 14872 2099 14875
rect 2222 14872 2228 14884
rect 2087 14844 2228 14872
rect 2087 14841 2099 14844
rect 2041 14835 2099 14841
rect 2222 14832 2228 14844
rect 2280 14832 2286 14884
rect 2133 14807 2191 14813
rect 2133 14773 2145 14807
rect 2179 14804 2191 14807
rect 2317 14807 2375 14813
rect 2317 14804 2329 14807
rect 2179 14776 2329 14804
rect 2179 14773 2191 14776
rect 2133 14767 2191 14773
rect 2317 14773 2329 14776
rect 2363 14804 2375 14807
rect 2746 14804 2774 14912
rect 2961 14909 2973 14912
rect 3007 14909 3019 14943
rect 2961 14903 3019 14909
rect 3602 14900 3608 14952
rect 3660 14900 3666 14952
rect 4157 14943 4215 14949
rect 4157 14909 4169 14943
rect 4203 14940 4215 14943
rect 4246 14940 4252 14952
rect 4203 14912 4252 14940
rect 4203 14909 4215 14912
rect 4157 14903 4215 14909
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 4341 14943 4399 14949
rect 4341 14909 4353 14943
rect 4387 14940 4399 14943
rect 4617 14943 4675 14949
rect 4387 14912 4476 14940
rect 4387 14909 4399 14912
rect 4341 14903 4399 14909
rect 2363 14776 2774 14804
rect 2363 14773 2375 14776
rect 2317 14767 2375 14773
rect 3050 14764 3056 14816
rect 3108 14764 3114 14816
rect 4062 14764 4068 14816
rect 4120 14764 4126 14816
rect 4448 14804 4476 14912
rect 4617 14909 4629 14943
rect 4663 14940 4675 14943
rect 4890 14940 4896 14952
rect 4663 14912 4896 14940
rect 4663 14909 4675 14912
rect 4617 14903 4675 14909
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5074 14900 5080 14952
rect 5132 14900 5138 14952
rect 6641 14943 6699 14949
rect 6641 14940 6653 14943
rect 6196 14912 6653 14940
rect 4522 14832 4528 14884
rect 4580 14872 4586 14884
rect 5258 14872 5264 14884
rect 4580 14844 5264 14872
rect 4580 14832 4586 14844
rect 5258 14832 5264 14844
rect 5316 14832 5322 14884
rect 6196 14881 6224 14912
rect 6641 14909 6653 14912
rect 6687 14909 6699 14943
rect 8389 14943 8447 14949
rect 8389 14940 8401 14943
rect 6641 14903 6699 14909
rect 7668 14912 8401 14940
rect 6181 14875 6239 14881
rect 6181 14841 6193 14875
rect 6227 14841 6239 14875
rect 6181 14835 6239 14841
rect 4614 14804 4620 14816
rect 4448 14776 4620 14804
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 4706 14764 4712 14816
rect 4764 14804 4770 14816
rect 4893 14807 4951 14813
rect 4893 14804 4905 14807
rect 4764 14776 4905 14804
rect 4764 14764 4770 14776
rect 4893 14773 4905 14776
rect 4939 14773 4951 14807
rect 4893 14767 4951 14773
rect 5997 14807 6055 14813
rect 5997 14773 6009 14807
rect 6043 14804 6055 14807
rect 6086 14804 6092 14816
rect 6043 14776 6092 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6086 14764 6092 14776
rect 6144 14764 6150 14816
rect 6362 14764 6368 14816
rect 6420 14804 6426 14816
rect 7668 14804 7696 14912
rect 8389 14909 8401 14912
rect 8435 14909 8447 14943
rect 9140 14940 9168 14971
rect 9582 14968 9588 15020
rect 9640 14968 9646 15020
rect 11716 15017 11744 15048
rect 11974 15036 11980 15088
rect 12032 15076 12038 15088
rect 12621 15079 12679 15085
rect 12621 15076 12633 15079
rect 12032 15048 12633 15076
rect 12032 15036 12038 15048
rect 12621 15045 12633 15048
rect 12667 15045 12679 15079
rect 12621 15039 12679 15045
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 12526 15008 12532 15020
rect 11747 14980 12532 15008
rect 11747 14977 11759 14980
rect 11701 14971 11759 14977
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 12728 15008 12756 15116
rect 13262 15104 13268 15156
rect 13320 15144 13326 15156
rect 13449 15147 13507 15153
rect 13449 15144 13461 15147
rect 13320 15116 13461 15144
rect 13320 15104 13326 15116
rect 13449 15113 13461 15116
rect 13495 15113 13507 15147
rect 13449 15107 13507 15113
rect 13538 15104 13544 15156
rect 13596 15144 13602 15156
rect 13596 15116 17540 15144
rect 13596 15104 13602 15116
rect 15470 15036 15476 15088
rect 15528 15076 15534 15088
rect 16025 15079 16083 15085
rect 16025 15076 16037 15079
rect 15528 15048 16037 15076
rect 15528 15036 15534 15048
rect 16025 15045 16037 15048
rect 16071 15045 16083 15079
rect 16025 15039 16083 15045
rect 16209 15079 16267 15085
rect 16209 15045 16221 15079
rect 16255 15076 16267 15079
rect 17402 15076 17408 15088
rect 16255 15048 17408 15076
rect 16255 15045 16267 15048
rect 16209 15039 16267 15045
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12728 14980 13001 15008
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 14977 13323 15011
rect 13265 14971 13323 14977
rect 9858 14940 9864 14952
rect 9140 14912 9864 14940
rect 8389 14903 8447 14909
rect 9858 14900 9864 14912
rect 9916 14940 9922 14952
rect 11054 14940 11060 14952
rect 9916 14912 11060 14940
rect 9916 14900 9922 14912
rect 11054 14900 11060 14912
rect 11112 14940 11118 14952
rect 11514 14940 11520 14952
rect 11112 14912 11520 14940
rect 11112 14900 11118 14912
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 11974 14900 11980 14952
rect 12032 14900 12038 14952
rect 12434 14900 12440 14952
rect 12492 14940 12498 14952
rect 13280 14940 13308 14971
rect 13538 14968 13544 15020
rect 13596 14968 13602 15020
rect 15197 15011 15255 15017
rect 15197 14977 15209 15011
rect 15243 15008 15255 15011
rect 15378 15008 15384 15020
rect 15243 14980 15384 15008
rect 15243 14977 15255 14980
rect 15197 14971 15255 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 12492 14912 13308 14940
rect 15565 14943 15623 14949
rect 12492 14900 12498 14912
rect 15565 14909 15577 14943
rect 15611 14940 15623 14943
rect 16224 14940 16252 15039
rect 16666 14968 16672 15020
rect 16724 14968 16730 15020
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 15008 17003 15011
rect 17034 15008 17040 15020
rect 16991 14980 17040 15008
rect 16991 14977 17003 14980
rect 16945 14971 17003 14977
rect 15611 14912 16252 14940
rect 16868 14940 16896 14971
rect 17034 14968 17040 14980
rect 17092 14968 17098 15020
rect 17144 15017 17172 15048
rect 17402 15036 17408 15048
rect 17460 15036 17466 15088
rect 17512 15076 17540 15116
rect 17586 15104 17592 15156
rect 17644 15104 17650 15156
rect 17681 15147 17739 15153
rect 17681 15113 17693 15147
rect 17727 15144 17739 15147
rect 17770 15144 17776 15156
rect 17727 15116 17776 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 17770 15104 17776 15116
rect 17828 15104 17834 15156
rect 17512 15048 18184 15076
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 17218 14968 17224 15020
rect 17276 14968 17282 15020
rect 17497 15011 17555 15017
rect 17497 14977 17509 15011
rect 17543 14977 17555 15011
rect 17497 14971 17555 14977
rect 17313 14943 17371 14949
rect 17313 14940 17325 14943
rect 16868 14912 17325 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 17313 14909 17325 14912
rect 17359 14909 17371 14943
rect 17313 14903 17371 14909
rect 9950 14832 9956 14884
rect 10008 14872 10014 14884
rect 10008 14844 12664 14872
rect 10008 14832 10014 14844
rect 6420 14776 7696 14804
rect 6420 14764 6426 14776
rect 8662 14764 8668 14816
rect 8720 14804 8726 14816
rect 9766 14804 9772 14816
rect 8720 14776 9772 14804
rect 8720 14764 8726 14776
rect 9766 14764 9772 14776
rect 9824 14804 9830 14816
rect 10226 14804 10232 14816
rect 9824 14776 10232 14804
rect 9824 14764 9830 14776
rect 10226 14764 10232 14776
rect 10284 14764 10290 14816
rect 12434 14764 12440 14816
rect 12492 14764 12498 14816
rect 12636 14813 12664 14844
rect 15470 14832 15476 14884
rect 15528 14832 15534 14884
rect 16666 14832 16672 14884
rect 16724 14872 16730 14884
rect 17512 14872 17540 14971
rect 18046 14968 18052 15020
rect 18104 15008 18110 15020
rect 18156 15017 18184 15048
rect 18141 15011 18199 15017
rect 18141 15008 18153 15011
rect 18104 14980 18153 15008
rect 18104 14968 18110 14980
rect 18141 14977 18153 14980
rect 18187 14977 18199 15011
rect 18141 14971 18199 14977
rect 18322 14968 18328 15020
rect 18380 14968 18386 15020
rect 18414 14968 18420 15020
rect 18472 14968 18478 15020
rect 16724 14844 17540 14872
rect 17865 14875 17923 14881
rect 16724 14832 16730 14844
rect 17865 14841 17877 14875
rect 17911 14872 17923 14875
rect 17954 14872 17960 14884
rect 17911 14844 17960 14872
rect 17911 14841 17923 14844
rect 17865 14835 17923 14841
rect 17954 14832 17960 14844
rect 18012 14832 18018 14884
rect 12621 14807 12679 14813
rect 12621 14773 12633 14807
rect 12667 14773 12679 14807
rect 12621 14767 12679 14773
rect 12802 14764 12808 14816
rect 12860 14804 12866 14816
rect 13173 14807 13231 14813
rect 13173 14804 13185 14807
rect 12860 14776 13185 14804
rect 12860 14764 12866 14776
rect 13173 14773 13185 14776
rect 13219 14773 13231 14807
rect 13173 14767 13231 14773
rect 15286 14764 15292 14816
rect 15344 14813 15350 14816
rect 15344 14807 15393 14813
rect 15344 14773 15347 14807
rect 15381 14773 15393 14807
rect 15344 14767 15393 14773
rect 15344 14764 15350 14767
rect 15838 14764 15844 14816
rect 15896 14764 15902 14816
rect 16390 14764 16396 14816
rect 16448 14764 16454 14816
rect 1104 14714 18860 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 18860 14714
rect 1104 14640 18860 14662
rect 2222 14560 2228 14612
rect 2280 14600 2286 14612
rect 2958 14600 2964 14612
rect 2280 14572 2964 14600
rect 2280 14560 2286 14572
rect 2958 14560 2964 14572
rect 3016 14600 3022 14612
rect 3878 14600 3884 14612
rect 3016 14572 3884 14600
rect 3016 14560 3022 14572
rect 3878 14560 3884 14572
rect 3936 14560 3942 14612
rect 3970 14560 3976 14612
rect 4028 14560 4034 14612
rect 4249 14603 4307 14609
rect 4249 14569 4261 14603
rect 4295 14600 4307 14603
rect 4614 14600 4620 14612
rect 4295 14572 4620 14600
rect 4295 14569 4307 14572
rect 4249 14563 4307 14569
rect 4614 14560 4620 14572
rect 4672 14560 4678 14612
rect 4798 14560 4804 14612
rect 4856 14560 4862 14612
rect 5074 14560 5080 14612
rect 5132 14560 5138 14612
rect 5994 14560 6000 14612
rect 6052 14560 6058 14612
rect 6288 14572 6684 14600
rect 1581 14535 1639 14541
rect 1581 14501 1593 14535
rect 1627 14532 1639 14535
rect 1670 14532 1676 14544
rect 1627 14504 1676 14532
rect 1627 14501 1639 14504
rect 1581 14495 1639 14501
rect 1670 14492 1676 14504
rect 1728 14532 1734 14544
rect 2038 14532 2044 14544
rect 1728 14504 2044 14532
rect 1728 14492 1734 14504
rect 2038 14492 2044 14504
rect 2096 14532 2102 14544
rect 2501 14535 2559 14541
rect 2501 14532 2513 14535
rect 2096 14504 2513 14532
rect 2096 14492 2102 14504
rect 2501 14501 2513 14504
rect 2547 14501 2559 14535
rect 3988 14532 4016 14560
rect 3988 14504 4200 14532
rect 2501 14495 2559 14501
rect 2222 14424 2228 14476
rect 2280 14424 2286 14476
rect 2685 14467 2743 14473
rect 2685 14433 2697 14467
rect 2731 14464 2743 14467
rect 3050 14464 3056 14476
rect 2731 14436 3056 14464
rect 2731 14433 2743 14436
rect 2685 14427 2743 14433
rect 3050 14424 3056 14436
rect 3108 14464 3114 14476
rect 3108 14436 4108 14464
rect 3108 14424 3114 14436
rect 842 14356 848 14408
rect 900 14396 906 14408
rect 1397 14399 1455 14405
rect 1397 14396 1409 14399
rect 900 14368 1409 14396
rect 900 14356 906 14368
rect 1397 14365 1409 14368
rect 1443 14365 1455 14399
rect 1397 14359 1455 14365
rect 3789 14399 3847 14405
rect 3789 14365 3801 14399
rect 3835 14396 3847 14399
rect 3878 14396 3884 14408
rect 3835 14368 3884 14396
rect 3835 14365 3847 14368
rect 3789 14359 3847 14365
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 4080 14405 4108 14436
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4065 14399 4123 14405
rect 4065 14365 4077 14399
rect 4111 14365 4123 14399
rect 4172 14396 4200 14504
rect 5810 14492 5816 14544
rect 5868 14532 5874 14544
rect 6288 14532 6316 14572
rect 5868 14504 6316 14532
rect 5868 14492 5874 14504
rect 6362 14492 6368 14544
rect 6420 14492 6426 14544
rect 6656 14532 6684 14572
rect 6730 14560 6736 14612
rect 6788 14560 6794 14612
rect 9950 14560 9956 14612
rect 10008 14560 10014 14612
rect 11903 14603 11961 14609
rect 11903 14569 11915 14603
rect 11949 14600 11961 14603
rect 12434 14600 12440 14612
rect 11949 14572 12440 14600
rect 11949 14569 11961 14572
rect 11903 14563 11961 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 13446 14560 13452 14612
rect 13504 14600 13510 14612
rect 15470 14600 15476 14612
rect 13504 14572 15476 14600
rect 13504 14560 13510 14572
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16485 14603 16543 14609
rect 16485 14600 16497 14603
rect 15804 14572 16497 14600
rect 15804 14560 15810 14572
rect 16485 14569 16497 14572
rect 16531 14569 16543 14603
rect 16485 14563 16543 14569
rect 16666 14560 16672 14612
rect 16724 14560 16730 14612
rect 17129 14603 17187 14609
rect 17129 14569 17141 14603
rect 17175 14600 17187 14603
rect 17218 14600 17224 14612
rect 17175 14572 17224 14600
rect 17175 14569 17187 14572
rect 17129 14563 17187 14569
rect 17218 14560 17224 14572
rect 17276 14560 17282 14612
rect 17313 14603 17371 14609
rect 17313 14569 17325 14603
rect 17359 14569 17371 14603
rect 17313 14563 17371 14569
rect 8662 14532 8668 14544
rect 6656 14504 8668 14532
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 12526 14492 12532 14544
rect 12584 14532 12590 14544
rect 17328 14532 17356 14563
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 17589 14603 17647 14609
rect 17589 14600 17601 14603
rect 17460 14572 17601 14600
rect 17460 14560 17466 14572
rect 17589 14569 17601 14572
rect 17635 14569 17647 14603
rect 17589 14563 17647 14569
rect 17773 14603 17831 14609
rect 17773 14569 17785 14603
rect 17819 14600 17831 14603
rect 18322 14600 18328 14612
rect 17819 14572 18328 14600
rect 17819 14569 17831 14572
rect 17773 14563 17831 14569
rect 18322 14560 18328 14572
rect 18380 14560 18386 14612
rect 17954 14532 17960 14544
rect 12584 14504 15240 14532
rect 12584 14492 12590 14504
rect 4433 14467 4491 14473
rect 4433 14433 4445 14467
rect 4479 14464 4491 14467
rect 4614 14464 4620 14476
rect 4479 14436 4620 14464
rect 4479 14433 4491 14436
rect 4433 14427 4491 14433
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 6380 14464 6408 14492
rect 6196 14436 6408 14464
rect 4249 14399 4307 14405
rect 4249 14396 4261 14399
rect 4172 14368 4261 14396
rect 4065 14359 4123 14365
rect 4249 14365 4261 14368
rect 4295 14365 4307 14399
rect 4249 14359 4307 14365
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 3602 14288 3608 14340
rect 3660 14328 3666 14340
rect 3988 14328 4016 14359
rect 3660 14300 4016 14328
rect 4540 14328 4568 14359
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 6196 14405 6224 14436
rect 10870 14424 10876 14476
rect 10928 14464 10934 14476
rect 12161 14467 12219 14473
rect 12161 14464 12173 14467
rect 10928 14436 12173 14464
rect 10928 14424 10934 14436
rect 12161 14433 12173 14436
rect 12207 14433 12219 14467
rect 13262 14464 13268 14476
rect 12161 14427 12219 14433
rect 13096 14436 13268 14464
rect 4893 14399 4951 14405
rect 4893 14396 4905 14399
rect 4856 14368 4905 14396
rect 4856 14356 4862 14368
rect 4893 14365 4905 14368
rect 4939 14365 4951 14399
rect 4893 14359 4951 14365
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14365 6239 14399
rect 6181 14359 6239 14365
rect 6270 14356 6276 14408
rect 6328 14396 6334 14408
rect 6365 14399 6423 14405
rect 6365 14396 6377 14399
rect 6328 14368 6377 14396
rect 6328 14356 6334 14368
rect 6365 14365 6377 14368
rect 6411 14365 6423 14399
rect 6365 14359 6423 14365
rect 13096 14392 13124 14436
rect 13262 14424 13268 14436
rect 13320 14424 13326 14476
rect 13354 14424 13360 14476
rect 13412 14464 13418 14476
rect 15212 14473 15240 14504
rect 15764 14504 16528 14532
rect 17328 14504 17960 14532
rect 15197 14467 15255 14473
rect 13412 14436 13952 14464
rect 13412 14424 13418 14436
rect 13173 14399 13231 14405
rect 13173 14392 13185 14399
rect 13096 14365 13185 14392
rect 13219 14365 13231 14399
rect 13446 14396 13452 14408
rect 13096 14364 13231 14365
rect 13173 14359 13231 14364
rect 13280 14368 13452 14396
rect 5442 14328 5448 14340
rect 4540 14300 5448 14328
rect 3660 14288 3666 14300
rect 3988 14272 4016 14300
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 8205 14331 8263 14337
rect 8205 14297 8217 14331
rect 8251 14328 8263 14331
rect 9582 14328 9588 14340
rect 8251 14300 9588 14328
rect 8251 14297 8263 14300
rect 8205 14291 8263 14297
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 10137 14331 10195 14337
rect 10137 14297 10149 14331
rect 10183 14297 10195 14331
rect 10137 14291 10195 14297
rect 3970 14220 3976 14272
rect 4028 14260 4034 14272
rect 5810 14260 5816 14272
rect 4028 14232 5816 14260
rect 4028 14220 4034 14232
rect 5810 14220 5816 14232
rect 5868 14220 5874 14272
rect 10152 14260 10180 14291
rect 10318 14288 10324 14340
rect 10376 14288 10382 14340
rect 12802 14328 12808 14340
rect 11454 14300 11560 14328
rect 10410 14260 10416 14272
rect 10152 14232 10416 14260
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 11532 14260 11560 14300
rect 11992 14300 12808 14328
rect 11992 14260 12020 14300
rect 12802 14288 12808 14300
rect 12860 14288 12866 14340
rect 13280 14337 13308 14368
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14398 13599 14399
rect 13648 14398 13676 14436
rect 13587 14370 13676 14398
rect 13817 14399 13875 14405
rect 13587 14365 13599 14370
rect 13541 14359 13599 14365
rect 13817 14365 13829 14399
rect 13863 14365 13875 14399
rect 13924 14396 13952 14436
rect 15197 14433 15209 14467
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 15764 14396 15792 14504
rect 15930 14424 15936 14476
rect 15988 14424 15994 14476
rect 16390 14424 16396 14476
rect 16448 14424 16454 14476
rect 16500 14464 16528 14504
rect 17954 14492 17960 14504
rect 18012 14492 18018 14544
rect 17770 14464 17776 14476
rect 16500 14436 17776 14464
rect 17770 14424 17776 14436
rect 17828 14424 17834 14476
rect 18414 14464 18420 14476
rect 17880 14436 18420 14464
rect 13924 14368 15792 14396
rect 13817 14359 13875 14365
rect 13265 14331 13323 14337
rect 12912 14300 13216 14328
rect 11532 14232 12020 14260
rect 12066 14220 12072 14272
rect 12124 14260 12130 14272
rect 12912 14260 12940 14300
rect 12124 14232 12940 14260
rect 12124 14220 12130 14232
rect 12986 14220 12992 14272
rect 13044 14220 13050 14272
rect 13188 14260 13216 14300
rect 13265 14297 13277 14331
rect 13311 14297 13323 14331
rect 13265 14291 13323 14297
rect 13357 14331 13415 14337
rect 13357 14297 13369 14331
rect 13403 14328 13415 14331
rect 13722 14328 13728 14340
rect 13403 14300 13728 14328
rect 13403 14297 13415 14300
rect 13357 14291 13415 14297
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 13832 14328 13860 14359
rect 15838 14356 15844 14408
rect 15896 14356 15902 14408
rect 16206 14356 16212 14408
rect 16264 14356 16270 14408
rect 17034 14356 17040 14408
rect 17092 14356 17098 14408
rect 17144 14368 17540 14396
rect 16574 14328 16580 14340
rect 13832 14300 16580 14328
rect 13832 14260 13860 14300
rect 16574 14288 16580 14300
rect 16632 14328 16638 14340
rect 17144 14328 17172 14368
rect 17310 14337 17316 14340
rect 16632 14300 17172 14328
rect 17297 14331 17316 14337
rect 16632 14288 16638 14300
rect 17297 14297 17309 14331
rect 17297 14291 17316 14297
rect 17310 14288 17316 14291
rect 17368 14288 17374 14340
rect 17512 14337 17540 14368
rect 17497 14331 17555 14337
rect 17497 14297 17509 14331
rect 17543 14297 17555 14331
rect 17497 14291 17555 14297
rect 17757 14331 17815 14337
rect 17757 14297 17769 14331
rect 17803 14328 17815 14331
rect 17880 14328 17908 14436
rect 18414 14424 18420 14436
rect 18472 14424 18478 14476
rect 18230 14356 18236 14408
rect 18288 14356 18294 14408
rect 18506 14356 18512 14408
rect 18564 14356 18570 14408
rect 17803 14300 17908 14328
rect 17803 14297 17815 14300
rect 17757 14291 17815 14297
rect 17954 14288 17960 14340
rect 18012 14288 18018 14340
rect 13188 14232 13860 14260
rect 16666 14220 16672 14272
rect 16724 14220 16730 14272
rect 17862 14220 17868 14272
rect 17920 14260 17926 14272
rect 18049 14263 18107 14269
rect 18049 14260 18061 14263
rect 17920 14232 18061 14260
rect 17920 14220 17926 14232
rect 18049 14229 18061 14232
rect 18095 14229 18107 14263
rect 18049 14223 18107 14229
rect 18325 14263 18383 14269
rect 18325 14229 18337 14263
rect 18371 14260 18383 14263
rect 18371 14232 18920 14260
rect 18371 14229 18383 14232
rect 18325 14223 18383 14229
rect 1104 14170 18860 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 18860 14170
rect 1104 14096 18860 14118
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 6362 14056 6368 14068
rect 5868 14028 6368 14056
rect 5868 14016 5874 14028
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 7650 14056 7656 14068
rect 7607 14028 7656 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 9858 14016 9864 14068
rect 9916 14056 9922 14068
rect 10163 14059 10221 14065
rect 10163 14056 10175 14059
rect 9916 14028 10175 14056
rect 9916 14016 9922 14028
rect 10163 14025 10175 14028
rect 10209 14056 10221 14059
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10209 14028 10609 14056
rect 10209 14025 10221 14028
rect 10163 14019 10221 14025
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 10597 14019 10655 14025
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 12338 14059 12396 14065
rect 10744 14028 12204 14056
rect 10744 14016 10750 14028
rect 6270 13988 6276 14000
rect 5736 13960 6276 13988
rect 5736 13932 5764 13960
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 6457 13991 6515 13997
rect 6457 13957 6469 13991
rect 6503 13988 6515 13991
rect 6730 13988 6736 14000
rect 6503 13960 6736 13988
rect 6503 13957 6515 13960
rect 6457 13951 6515 13957
rect 6730 13948 6736 13960
rect 6788 13948 6794 14000
rect 8662 13948 8668 14000
rect 8720 13988 8726 14000
rect 8941 13991 8999 13997
rect 8941 13988 8953 13991
rect 8720 13960 8953 13988
rect 8720 13948 8726 13960
rect 8941 13957 8953 13960
rect 8987 13957 8999 13991
rect 8941 13951 8999 13957
rect 9122 13948 9128 14000
rect 9180 13997 9186 14000
rect 9180 13991 9199 13997
rect 9187 13957 9199 13991
rect 9180 13951 9199 13957
rect 9953 13991 10011 13997
rect 9953 13957 9965 13991
rect 9999 13957 10011 13991
rect 9953 13951 10011 13957
rect 9180 13948 9186 13951
rect 2038 13880 2044 13932
rect 2096 13880 2102 13932
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 2225 13923 2283 13929
rect 2225 13920 2237 13923
rect 2188 13892 2237 13920
rect 2188 13880 2194 13892
rect 2225 13889 2237 13892
rect 2271 13920 2283 13923
rect 2590 13920 2596 13932
rect 2271 13892 2596 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 5718 13880 5724 13932
rect 5776 13880 5782 13932
rect 5997 13923 6055 13929
rect 5997 13889 6009 13923
rect 6043 13920 6055 13923
rect 6546 13920 6552 13932
rect 6043 13892 6552 13920
rect 6043 13889 6055 13892
rect 5997 13883 6055 13889
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13920 7711 13923
rect 7742 13920 7748 13932
rect 7699 13892 7748 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 9968 13852 9996 13951
rect 10410 13948 10416 14000
rect 10468 13988 10474 14000
rect 10965 13991 11023 13997
rect 10965 13988 10977 13991
rect 10468 13960 10977 13988
rect 10468 13948 10474 13960
rect 10965 13957 10977 13960
rect 11011 13988 11023 13991
rect 12066 13988 12072 14000
rect 11011 13960 12072 13988
rect 11011 13957 11023 13960
rect 10965 13951 11023 13957
rect 12066 13948 12072 13960
rect 12124 13948 12130 14000
rect 12176 13929 12204 14028
rect 12338 14025 12350 14059
rect 12384 14056 12396 14059
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12384 14028 12909 14056
rect 12384 14025 12396 14028
rect 12338 14019 12396 14025
rect 12897 14025 12909 14028
rect 12943 14025 12955 14059
rect 12897 14019 12955 14025
rect 15473 14059 15531 14065
rect 15473 14025 15485 14059
rect 15519 14056 15531 14059
rect 16666 14056 16672 14068
rect 15519 14028 16672 14056
rect 15519 14025 15531 14028
rect 15473 14019 15531 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17037 14059 17095 14065
rect 17037 14056 17049 14059
rect 16816 14028 17049 14056
rect 16816 14016 16822 14028
rect 17037 14025 17049 14028
rect 17083 14025 17095 14059
rect 17037 14019 17095 14025
rect 18049 14059 18107 14065
rect 18049 14025 18061 14059
rect 18095 14056 18107 14059
rect 18322 14056 18328 14068
rect 18095 14028 18328 14056
rect 18095 14025 18107 14028
rect 18049 14019 18107 14025
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 18414 14016 18420 14068
rect 18472 14016 18478 14068
rect 12437 13991 12495 13997
rect 12437 13957 12449 13991
rect 12483 13988 12495 13991
rect 12618 13988 12624 14000
rect 12483 13960 12624 13988
rect 12483 13957 12495 13960
rect 12437 13951 12495 13957
rect 12618 13948 12624 13960
rect 12676 13988 12682 14000
rect 12986 13988 12992 14000
rect 12676 13960 12992 13988
rect 12676 13948 12682 13960
rect 12986 13948 12992 13960
rect 13044 13948 13050 14000
rect 13081 13991 13139 13997
rect 13081 13957 13093 13991
rect 13127 13988 13139 13991
rect 13170 13988 13176 14000
rect 13127 13960 13176 13988
rect 13127 13957 13139 13960
rect 13081 13951 13139 13957
rect 13170 13948 13176 13960
rect 13228 13948 13234 14000
rect 14001 13991 14059 13997
rect 14001 13988 14013 13991
rect 13280 13960 14013 13988
rect 10781 13923 10839 13929
rect 10781 13889 10793 13923
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13889 12219 13923
rect 12161 13883 12219 13889
rect 12253 13923 12311 13929
rect 12253 13889 12265 13923
rect 12299 13920 12311 13923
rect 12713 13923 12771 13929
rect 12299 13892 12434 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 10502 13852 10508 13864
rect 9968 13824 10508 13852
rect 10502 13812 10508 13824
rect 10560 13852 10566 13864
rect 10796 13852 10824 13883
rect 12066 13852 12072 13864
rect 10560 13824 12072 13852
rect 10560 13812 10566 13824
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 10686 13784 10692 13796
rect 10152 13756 10692 13784
rect 10152 13728 10180 13756
rect 10686 13744 10692 13756
rect 10744 13744 10750 13796
rect 12176 13784 12204 13883
rect 12406 13864 12434 13892
rect 12713 13889 12725 13923
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 12406 13824 12440 13864
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 12526 13812 12532 13864
rect 12584 13812 12590 13864
rect 12728 13852 12756 13883
rect 12802 13880 12808 13932
rect 12860 13880 12866 13932
rect 13280 13852 13308 13960
rect 14001 13957 14013 13960
rect 14047 13957 14059 13991
rect 15749 13991 15807 13997
rect 15749 13988 15761 13991
rect 14001 13951 14059 13957
rect 15120 13960 15761 13988
rect 15120 13932 15148 13960
rect 15749 13957 15761 13960
rect 15795 13957 15807 13991
rect 15749 13951 15807 13957
rect 15841 13991 15899 13997
rect 15841 13957 15853 13991
rect 15887 13988 15899 13991
rect 16853 13991 16911 13997
rect 16853 13988 16865 13991
rect 15887 13960 16865 13988
rect 15887 13957 15899 13960
rect 15841 13951 15899 13957
rect 16853 13957 16865 13960
rect 16899 13957 16911 13991
rect 16853 13951 16911 13957
rect 17604 13960 17908 13988
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 13446 13880 13452 13932
rect 13504 13880 13510 13932
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 13556 13892 13921 13920
rect 12728 13824 13308 13852
rect 13078 13784 13084 13796
rect 12176 13756 13084 13784
rect 13078 13744 13084 13756
rect 13136 13744 13142 13796
rect 13173 13787 13231 13793
rect 13173 13753 13185 13787
rect 13219 13784 13231 13787
rect 13556 13784 13584 13892
rect 13909 13889 13921 13892
rect 13955 13889 13967 13923
rect 13909 13883 13967 13889
rect 15102 13880 15108 13932
rect 15160 13880 15166 13932
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 15252 13892 15301 13920
rect 15252 13880 15258 13892
rect 15289 13889 15301 13892
rect 15335 13920 15347 13923
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 15335 13892 15577 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 15565 13889 15577 13892
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 13725 13855 13783 13861
rect 13725 13821 13737 13855
rect 13771 13821 13783 13855
rect 13725 13815 13783 13821
rect 13219 13756 13584 13784
rect 13740 13784 13768 13815
rect 13814 13812 13820 13864
rect 13872 13852 13878 13864
rect 15856 13852 15884 13951
rect 15933 13923 15991 13929
rect 15933 13889 15945 13923
rect 15979 13920 15991 13923
rect 16114 13920 16120 13932
rect 15979 13892 16120 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16114 13880 16120 13892
rect 16172 13920 16178 13932
rect 17604 13929 17632 13960
rect 17880 13932 17908 13960
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16172 13892 16681 13920
rect 16172 13880 16178 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 17034 13852 17040 13864
rect 13872 13824 15884 13852
rect 16132 13824 17040 13852
rect 13872 13812 13878 13824
rect 16132 13793 16160 13824
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17696 13796 17724 13883
rect 17862 13880 17868 13932
rect 17920 13920 17926 13932
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 17920 13892 18153 13920
rect 17920 13880 17926 13892
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 17770 13812 17776 13864
rect 17828 13852 17834 13864
rect 18417 13855 18475 13861
rect 18417 13852 18429 13855
rect 17828 13824 18429 13852
rect 17828 13812 17834 13824
rect 18417 13821 18429 13824
rect 18463 13852 18475 13855
rect 18892 13852 18920 14232
rect 18463 13824 18920 13852
rect 18463 13821 18475 13824
rect 18417 13815 18475 13821
rect 16117 13787 16175 13793
rect 13740 13756 13860 13784
rect 13219 13753 13231 13756
rect 13173 13747 13231 13753
rect 2133 13719 2191 13725
rect 2133 13685 2145 13719
rect 2179 13716 2191 13719
rect 2590 13716 2596 13728
rect 2179 13688 2596 13716
rect 2179 13685 2191 13688
rect 2133 13679 2191 13685
rect 2590 13676 2596 13688
rect 2648 13676 2654 13728
rect 6181 13719 6239 13725
rect 6181 13685 6193 13719
rect 6227 13716 6239 13719
rect 6362 13716 6368 13728
rect 6227 13688 6368 13716
rect 6227 13685 6239 13688
rect 6181 13679 6239 13685
rect 6362 13676 6368 13688
rect 6420 13676 6426 13728
rect 8662 13676 8668 13728
rect 8720 13716 8726 13728
rect 9125 13719 9183 13725
rect 9125 13716 9137 13719
rect 8720 13688 9137 13716
rect 8720 13676 8726 13688
rect 9125 13685 9137 13688
rect 9171 13685 9183 13719
rect 9125 13679 9183 13685
rect 9214 13676 9220 13728
rect 9272 13716 9278 13728
rect 9309 13719 9367 13725
rect 9309 13716 9321 13719
rect 9272 13688 9321 13716
rect 9272 13676 9278 13688
rect 9309 13685 9321 13688
rect 9355 13685 9367 13719
rect 9309 13679 9367 13685
rect 10134 13676 10140 13728
rect 10192 13676 10198 13728
rect 10318 13676 10324 13728
rect 10376 13676 10382 13728
rect 10413 13719 10471 13725
rect 10413 13685 10425 13719
rect 10459 13716 10471 13719
rect 10962 13716 10968 13728
rect 10459 13688 10968 13716
rect 10459 13685 10471 13688
rect 10413 13679 10471 13685
rect 10962 13676 10968 13688
rect 11020 13676 11026 13728
rect 12986 13676 12992 13728
rect 13044 13716 13050 13728
rect 13188 13716 13216 13747
rect 13832 13728 13860 13756
rect 16117 13753 16129 13787
rect 16163 13753 16175 13787
rect 16117 13747 16175 13753
rect 17678 13744 17684 13796
rect 17736 13784 17742 13796
rect 18233 13787 18291 13793
rect 18233 13784 18245 13787
rect 17736 13756 18245 13784
rect 17736 13744 17742 13756
rect 18233 13753 18245 13756
rect 18279 13753 18291 13787
rect 18233 13747 18291 13753
rect 13044 13688 13216 13716
rect 13044 13676 13050 13688
rect 13814 13676 13820 13728
rect 13872 13676 13878 13728
rect 17494 13676 17500 13728
rect 17552 13676 17558 13728
rect 17862 13676 17868 13728
rect 17920 13676 17926 13728
rect 1104 13626 18860 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 18860 13626
rect 1104 13552 18860 13574
rect 4433 13515 4491 13521
rect 4433 13481 4445 13515
rect 4479 13512 4491 13515
rect 4798 13512 4804 13524
rect 4479 13484 4804 13512
rect 4479 13481 4491 13484
rect 4433 13475 4491 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5721 13515 5779 13521
rect 5721 13481 5733 13515
rect 5767 13512 5779 13515
rect 5810 13512 5816 13524
rect 5767 13484 5816 13512
rect 5767 13481 5779 13484
rect 5721 13475 5779 13481
rect 5810 13472 5816 13484
rect 5868 13472 5874 13524
rect 6362 13472 6368 13524
rect 6420 13472 6426 13524
rect 6546 13472 6552 13524
rect 6604 13512 6610 13524
rect 8389 13515 8447 13521
rect 8389 13512 8401 13515
rect 6604 13484 8401 13512
rect 6604 13472 6610 13484
rect 8389 13481 8401 13484
rect 8435 13481 8447 13515
rect 8389 13475 8447 13481
rect 8662 13472 8668 13524
rect 8720 13472 8726 13524
rect 10686 13512 10692 13524
rect 8864 13484 10692 13512
rect 2590 13404 2596 13456
rect 2648 13404 2654 13456
rect 3326 13404 3332 13456
rect 3384 13444 3390 13456
rect 3384 13416 4016 13444
rect 3384 13404 3390 13416
rect 3988 13388 4016 13416
rect 2038 13376 2044 13388
rect 1964 13348 2044 13376
rect 1394 13268 1400 13320
rect 1452 13268 1458 13320
rect 1964 13317 1992 13348
rect 2038 13336 2044 13348
rect 2096 13376 2102 13388
rect 2682 13376 2688 13388
rect 2096 13348 2688 13376
rect 2096 13336 2102 13348
rect 2682 13336 2688 13348
rect 2740 13336 2746 13388
rect 2777 13379 2835 13385
rect 2777 13345 2789 13379
rect 2823 13376 2835 13379
rect 2823 13348 3464 13376
rect 2823 13345 2835 13348
rect 2777 13339 2835 13345
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 2130 13268 2136 13320
rect 2188 13268 2194 13320
rect 3050 13268 3056 13320
rect 3108 13268 3114 13320
rect 3326 13268 3332 13320
rect 3384 13268 3390 13320
rect 3436 13317 3464 13348
rect 3970 13336 3976 13388
rect 4028 13376 4034 13388
rect 6564 13376 6592 13472
rect 4028 13348 4108 13376
rect 4028 13336 4034 13348
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 3510 13308 3516 13320
rect 3467 13280 3516 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 3878 13268 3884 13320
rect 3936 13268 3942 13320
rect 2317 13243 2375 13249
rect 2317 13240 2329 13243
rect 2240 13212 2329 13240
rect 2240 13184 2268 13212
rect 2317 13209 2329 13212
rect 2363 13209 2375 13243
rect 2317 13203 2375 13209
rect 3234 13200 3240 13252
rect 3292 13200 3298 13252
rect 4080 13249 4108 13348
rect 5552 13348 6592 13376
rect 4249 13311 4307 13317
rect 4249 13277 4261 13311
rect 4295 13308 4307 13311
rect 5552 13308 5580 13348
rect 6638 13336 6644 13388
rect 6696 13336 6702 13388
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 4295 13280 5580 13308
rect 4295 13277 4307 13280
rect 4249 13271 4307 13277
rect 4065 13243 4123 13249
rect 4065 13209 4077 13243
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4154 13200 4160 13252
rect 4212 13200 4218 13252
rect 5552 13249 5580 13280
rect 5920 13280 6009 13308
rect 5537 13243 5595 13249
rect 5537 13209 5549 13243
rect 5583 13240 5595 13243
rect 5626 13240 5632 13252
rect 5583 13212 5632 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 5626 13200 5632 13212
rect 5684 13200 5690 13252
rect 5718 13200 5724 13252
rect 5776 13249 5782 13252
rect 5776 13243 5795 13249
rect 5783 13209 5795 13243
rect 5776 13203 5795 13209
rect 5776 13200 5782 13203
rect 5920 13184 5948 13280
rect 5997 13277 6009 13280
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13277 8631 13311
rect 8573 13271 8631 13277
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 8864 13308 8892 13484
rect 10686 13472 10692 13484
rect 10744 13472 10750 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13265 13515 13323 13521
rect 13265 13512 13277 13515
rect 12860 13484 13277 13512
rect 12860 13472 12866 13484
rect 12710 13404 12716 13456
rect 12768 13444 12774 13456
rect 12989 13447 13047 13453
rect 12989 13444 13001 13447
rect 12768 13416 13001 13444
rect 12768 13404 12774 13416
rect 12989 13413 13001 13416
rect 13035 13413 13047 13447
rect 12989 13407 13047 13413
rect 8941 13379 8999 13385
rect 8941 13345 8953 13379
rect 8987 13376 8999 13379
rect 10870 13376 10876 13388
rect 8987 13348 10876 13376
rect 8987 13345 8999 13348
rect 8941 13339 8999 13345
rect 10870 13336 10876 13348
rect 10928 13336 10934 13388
rect 8803 13280 8892 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 6917 13243 6975 13249
rect 6917 13209 6929 13243
rect 6963 13209 6975 13243
rect 6917 13203 6975 13209
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 900 13144 1593 13172
rect 900 13132 906 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 2041 13175 2099 13181
rect 2041 13141 2053 13175
rect 2087 13172 2099 13175
rect 2222 13172 2228 13184
rect 2087 13144 2228 13172
rect 2087 13141 2099 13144
rect 2041 13135 2099 13141
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 3605 13175 3663 13181
rect 3605 13141 3617 13175
rect 3651 13172 3663 13175
rect 3970 13172 3976 13184
rect 3651 13144 3976 13172
rect 3651 13141 3663 13144
rect 3605 13135 3663 13141
rect 3970 13132 3976 13144
rect 4028 13132 4034 13184
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 6362 13132 6368 13184
rect 6420 13132 6426 13184
rect 6549 13175 6607 13181
rect 6549 13141 6561 13175
rect 6595 13172 6607 13175
rect 6932 13172 6960 13203
rect 7926 13200 7932 13252
rect 7984 13200 7990 13252
rect 6595 13144 6960 13172
rect 8588 13172 8616 13271
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12676 13280 12725 13308
rect 12676 13268 12682 13280
rect 12713 13277 12725 13280
rect 12759 13277 12771 13311
rect 12713 13271 12771 13277
rect 12986 13268 12992 13320
rect 13044 13268 13050 13320
rect 13188 13317 13216 13484
rect 13265 13481 13277 13484
rect 13311 13481 13323 13515
rect 13265 13475 13323 13481
rect 13722 13472 13728 13524
rect 13780 13472 13786 13524
rect 17129 13515 17187 13521
rect 17129 13481 17141 13515
rect 17175 13512 17187 13515
rect 17310 13512 17316 13524
rect 17175 13484 17316 13512
rect 17175 13481 17187 13484
rect 17129 13475 17187 13481
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 16574 13336 16580 13388
rect 16632 13376 16638 13388
rect 17313 13379 17371 13385
rect 17313 13376 17325 13379
rect 16632 13348 17325 13376
rect 16632 13336 16638 13348
rect 17313 13345 17325 13348
rect 17359 13376 17371 13379
rect 17678 13376 17684 13388
rect 17359 13348 17684 13376
rect 17359 13345 17371 13348
rect 17313 13339 17371 13345
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13277 13231 13311
rect 13173 13271 13231 13277
rect 13449 13311 13507 13317
rect 13449 13277 13461 13311
rect 13495 13277 13507 13311
rect 13449 13271 13507 13277
rect 9214 13200 9220 13252
rect 9272 13200 9278 13252
rect 9766 13200 9772 13252
rect 9824 13200 9830 13252
rect 11146 13200 11152 13252
rect 11204 13200 11210 13252
rect 11790 13200 11796 13252
rect 11848 13200 11854 13252
rect 13078 13200 13084 13252
rect 13136 13240 13142 13252
rect 13464 13240 13492 13271
rect 13538 13268 13544 13320
rect 13596 13268 13602 13320
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 17405 13311 17463 13317
rect 17405 13308 17417 13311
rect 13872 13280 17417 13308
rect 13872 13268 13878 13280
rect 17405 13277 17417 13280
rect 17451 13308 17463 13311
rect 17494 13308 17500 13320
rect 17451 13280 17500 13308
rect 17451 13277 17463 13280
rect 17405 13271 17463 13277
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 18506 13268 18512 13320
rect 18564 13268 18570 13320
rect 15194 13240 15200 13252
rect 13136 13212 15200 13240
rect 13136 13200 13142 13212
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 9858 13172 9864 13184
rect 8588 13144 9864 13172
rect 6595 13141 6607 13144
rect 6549 13135 6607 13141
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12621 13175 12679 13181
rect 12621 13172 12633 13175
rect 12124 13144 12633 13172
rect 12124 13132 12130 13144
rect 12621 13141 12633 13144
rect 12667 13172 12679 13175
rect 13722 13172 13728 13184
rect 12667 13144 13728 13172
rect 12667 13141 12679 13144
rect 12621 13135 12679 13141
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 18325 13175 18383 13181
rect 18325 13141 18337 13175
rect 18371 13172 18383 13175
rect 18414 13172 18420 13184
rect 18371 13144 18420 13172
rect 18371 13141 18383 13144
rect 18325 13135 18383 13141
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 1104 13082 18860 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 18860 13082
rect 1104 13008 18860 13030
rect 2409 12971 2467 12977
rect 2409 12937 2421 12971
rect 2455 12968 2467 12971
rect 3234 12968 3240 12980
rect 2455 12940 3240 12968
rect 2455 12937 2467 12940
rect 2409 12931 2467 12937
rect 3234 12928 3240 12940
rect 3292 12968 3298 12980
rect 3292 12940 4200 12968
rect 3292 12928 3298 12940
rect 2056 12872 2912 12900
rect 2056 12844 2084 12872
rect 1581 12835 1639 12841
rect 1581 12801 1593 12835
rect 1627 12801 1639 12835
rect 1581 12795 1639 12801
rect 1596 12708 1624 12795
rect 2038 12792 2044 12844
rect 2096 12792 2102 12844
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12801 2559 12835
rect 2501 12795 2559 12801
rect 2884 12832 2912 12872
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 2884 12804 3341 12832
rect 2133 12767 2191 12773
rect 2133 12733 2145 12767
rect 2179 12764 2191 12767
rect 2222 12764 2228 12776
rect 2179 12736 2228 12764
rect 2179 12733 2191 12736
rect 2133 12727 2191 12733
rect 2222 12724 2228 12736
rect 2280 12724 2286 12776
rect 1578 12656 1584 12708
rect 1636 12696 1642 12708
rect 2516 12696 2544 12795
rect 2682 12724 2688 12776
rect 2740 12764 2746 12776
rect 2884 12773 2912 12804
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 3786 12792 3792 12844
rect 3844 12792 3850 12844
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 4062 12792 4068 12844
rect 4120 12792 4126 12844
rect 4172 12841 4200 12940
rect 4614 12928 4620 12980
rect 4672 12928 4678 12980
rect 5626 12928 5632 12980
rect 5684 12928 5690 12980
rect 5718 12928 5724 12980
rect 5776 12968 5782 12980
rect 5813 12971 5871 12977
rect 5813 12968 5825 12971
rect 5776 12940 5825 12968
rect 5776 12928 5782 12940
rect 5813 12937 5825 12940
rect 5859 12937 5871 12971
rect 5813 12931 5871 12937
rect 5902 12928 5908 12980
rect 5960 12968 5966 12980
rect 7837 12971 7895 12977
rect 5960 12940 7052 12968
rect 5960 12928 5966 12940
rect 5644 12900 5672 12928
rect 4356 12872 5672 12900
rect 4356 12841 4384 12872
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12801 4399 12835
rect 4341 12795 4399 12801
rect 2869 12767 2927 12773
rect 2740 12736 2820 12764
rect 2740 12724 2746 12736
rect 2792 12705 2820 12736
rect 2869 12733 2881 12767
rect 2915 12733 2927 12767
rect 2869 12727 2927 12733
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3421 12767 3479 12773
rect 3421 12764 3433 12767
rect 3016 12736 3433 12764
rect 3016 12724 3022 12736
rect 3421 12733 3433 12736
rect 3467 12764 3479 12767
rect 3878 12764 3884 12776
rect 3467 12736 3884 12764
rect 3467 12733 3479 12736
rect 3421 12727 3479 12733
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 4356 12764 4384 12795
rect 4706 12792 4712 12844
rect 4764 12832 4770 12844
rect 5184 12841 5212 12872
rect 6362 12860 6368 12912
rect 6420 12900 6426 12912
rect 7024 12909 7052 12940
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 7926 12968 7932 12980
rect 7883 12940 7932 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 7926 12928 7932 12940
rect 7984 12928 7990 12980
rect 9122 12928 9128 12980
rect 9180 12968 9186 12980
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 9180 12940 9229 12968
rect 9180 12928 9186 12940
rect 9217 12937 9229 12940
rect 9263 12937 9275 12971
rect 9674 12968 9680 12980
rect 9217 12931 9275 12937
rect 9324 12940 9680 12968
rect 6733 12903 6791 12909
rect 6733 12900 6745 12903
rect 6420 12872 6745 12900
rect 6420 12860 6426 12872
rect 6733 12869 6745 12872
rect 6779 12869 6791 12903
rect 6733 12863 6791 12869
rect 7009 12903 7067 12909
rect 7009 12869 7021 12903
rect 7055 12869 7067 12903
rect 9324 12900 9352 12940
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 9766 12928 9772 12980
rect 9824 12928 9830 12980
rect 10873 12971 10931 12977
rect 10873 12937 10885 12971
rect 10919 12968 10931 12971
rect 11146 12968 11152 12980
rect 10919 12940 11152 12968
rect 10919 12937 10931 12940
rect 10873 12931 10931 12937
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11790 12928 11796 12980
rect 11848 12928 11854 12980
rect 12434 12928 12440 12980
rect 12492 12968 12498 12980
rect 13538 12968 13544 12980
rect 12492 12940 13544 12968
rect 12492 12928 12498 12940
rect 13538 12928 13544 12940
rect 13596 12968 13602 12980
rect 14093 12971 14151 12977
rect 14093 12968 14105 12971
rect 13596 12940 14105 12968
rect 13596 12928 13602 12940
rect 14093 12937 14105 12940
rect 14139 12968 14151 12971
rect 15654 12968 15660 12980
rect 14139 12940 15660 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 15654 12928 15660 12940
rect 15712 12928 15718 12980
rect 16114 12928 16120 12980
rect 16172 12928 16178 12980
rect 16574 12928 16580 12980
rect 16632 12968 16638 12980
rect 18049 12971 18107 12977
rect 18049 12968 18061 12971
rect 16632 12940 18061 12968
rect 16632 12928 16638 12940
rect 18049 12937 18061 12940
rect 18095 12937 18107 12971
rect 18049 12931 18107 12937
rect 7009 12863 7067 12869
rect 7116 12872 9352 12900
rect 9585 12903 9643 12909
rect 4801 12835 4859 12841
rect 4801 12832 4813 12835
rect 4764 12804 4813 12832
rect 4764 12792 4770 12804
rect 4801 12801 4813 12804
rect 4847 12801 4859 12835
rect 5077 12835 5135 12841
rect 5077 12832 5089 12835
rect 4801 12795 4859 12801
rect 4908 12804 5089 12832
rect 3988 12736 4384 12764
rect 4525 12767 4583 12773
rect 3988 12708 4016 12736
rect 4525 12733 4537 12767
rect 4571 12764 4583 12767
rect 4614 12764 4620 12776
rect 4571 12736 4620 12764
rect 4571 12733 4583 12736
rect 4525 12727 4583 12733
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 4908 12764 4936 12804
rect 5077 12801 5089 12804
rect 5123 12801 5135 12835
rect 5077 12795 5135 12801
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12801 5227 12835
rect 5169 12795 5227 12801
rect 5353 12835 5411 12841
rect 5353 12801 5365 12835
rect 5399 12832 5411 12835
rect 5534 12832 5540 12844
rect 5399 12804 5540 12832
rect 5399 12801 5411 12804
rect 5353 12795 5411 12801
rect 5534 12792 5540 12804
rect 5592 12792 5598 12844
rect 5721 12835 5779 12841
rect 5721 12801 5733 12835
rect 5767 12832 5779 12835
rect 5810 12832 5816 12844
rect 5767 12804 5816 12832
rect 5767 12801 5779 12804
rect 5721 12795 5779 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 6748 12832 6776 12863
rect 7116 12832 7144 12872
rect 9585 12869 9597 12903
rect 9631 12900 9643 12903
rect 9858 12900 9864 12912
rect 9631 12872 9864 12900
rect 9631 12869 9643 12872
rect 9585 12863 9643 12869
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 10686 12860 10692 12912
rect 10744 12860 10750 12912
rect 13998 12860 14004 12912
rect 14056 12900 14062 12912
rect 14210 12903 14268 12909
rect 14210 12900 14222 12903
rect 14056 12872 14222 12900
rect 14056 12860 14062 12872
rect 14210 12869 14222 12872
rect 14256 12900 14268 12903
rect 15010 12900 15016 12912
rect 14256 12872 15016 12900
rect 14256 12869 14268 12872
rect 14210 12863 14268 12869
rect 15010 12860 15016 12872
rect 15068 12860 15074 12912
rect 17494 12900 17500 12912
rect 15120 12872 17500 12900
rect 6748 12804 7144 12832
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 7742 12792 7748 12844
rect 7800 12832 7806 12844
rect 7926 12832 7932 12844
rect 7800 12804 7932 12832
rect 7800 12792 7806 12804
rect 7926 12792 7932 12804
rect 7984 12792 7990 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12801 9459 12835
rect 9401 12795 9459 12801
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12832 9735 12835
rect 9723 12804 10272 12832
rect 9723 12801 9735 12804
rect 9677 12795 9735 12801
rect 4724 12736 4936 12764
rect 1636 12668 2544 12696
rect 2777 12699 2835 12705
rect 1636 12656 1642 12668
rect 2777 12665 2789 12699
rect 2823 12665 2835 12699
rect 2777 12659 2835 12665
rect 3050 12656 3056 12708
rect 3108 12696 3114 12708
rect 3970 12696 3976 12708
rect 3108 12668 3976 12696
rect 3108 12656 3114 12668
rect 3970 12656 3976 12668
rect 4028 12656 4034 12708
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 4724 12696 4752 12736
rect 4982 12724 4988 12776
rect 5040 12764 5046 12776
rect 5445 12767 5503 12773
rect 5445 12764 5457 12767
rect 5040 12736 5457 12764
rect 5040 12724 5046 12736
rect 5445 12733 5457 12736
rect 5491 12764 5503 12767
rect 7208 12764 7236 12792
rect 5491 12736 7236 12764
rect 9416 12764 9444 12795
rect 10134 12764 10140 12776
rect 9416 12736 10140 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 10134 12724 10140 12736
rect 10192 12724 10198 12776
rect 10244 12764 10272 12804
rect 10318 12792 10324 12844
rect 10376 12792 10382 12844
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 11054 12764 11060 12776
rect 10244 12736 11060 12764
rect 11054 12724 11060 12736
rect 11112 12764 11118 12776
rect 11716 12764 11744 12795
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13412 12804 13737 12832
rect 13412 12792 13418 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 15120 12832 15148 12872
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 18325 12903 18383 12909
rect 18325 12900 18337 12903
rect 17604 12872 18337 12900
rect 13725 12795 13783 12801
rect 14768 12804 15148 12832
rect 11112 12736 11744 12764
rect 11112 12724 11118 12736
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14001 12767 14059 12773
rect 14001 12764 14013 12767
rect 13872 12736 14013 12764
rect 13872 12724 13878 12736
rect 14001 12733 14013 12736
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 4120 12668 4752 12696
rect 6365 12699 6423 12705
rect 4120 12656 4126 12668
rect 6365 12665 6377 12699
rect 6411 12665 6423 12699
rect 7377 12699 7435 12705
rect 7377 12696 7389 12699
rect 6365 12659 6423 12665
rect 6748 12668 7389 12696
rect 1670 12588 1676 12640
rect 1728 12588 1734 12640
rect 2130 12588 2136 12640
rect 2188 12628 2194 12640
rect 2639 12631 2697 12637
rect 2639 12628 2651 12631
rect 2188 12600 2651 12628
rect 2188 12588 2194 12600
rect 2639 12597 2651 12600
rect 2685 12597 2697 12631
rect 2639 12591 2697 12597
rect 2866 12588 2872 12640
rect 2924 12628 2930 12640
rect 2961 12631 3019 12637
rect 2961 12628 2973 12631
rect 2924 12600 2973 12628
rect 2924 12588 2930 12600
rect 2961 12597 2973 12600
rect 3007 12597 3019 12631
rect 2961 12591 3019 12597
rect 5902 12588 5908 12640
rect 5960 12628 5966 12640
rect 5997 12631 6055 12637
rect 5997 12628 6009 12631
rect 5960 12600 6009 12628
rect 5960 12588 5966 12600
rect 5997 12597 6009 12600
rect 6043 12628 6055 12631
rect 6380 12628 6408 12659
rect 6748 12637 6776 12668
rect 7377 12665 7389 12668
rect 7423 12665 7435 12699
rect 7377 12659 7435 12665
rect 14369 12699 14427 12705
rect 14369 12665 14381 12699
rect 14415 12696 14427 12699
rect 14461 12699 14519 12705
rect 14461 12696 14473 12699
rect 14415 12668 14473 12696
rect 14415 12665 14427 12668
rect 14369 12659 14427 12665
rect 14461 12665 14473 12668
rect 14507 12696 14519 12699
rect 14642 12696 14648 12708
rect 14507 12668 14648 12696
rect 14507 12665 14519 12668
rect 14461 12659 14519 12665
rect 14642 12656 14648 12668
rect 14700 12656 14706 12708
rect 14768 12696 14796 12804
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12832 16359 12835
rect 16347 12804 16712 12832
rect 16347 12801 16359 12804
rect 16301 12795 16359 12801
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 15488 12764 15516 12792
rect 15059 12736 15516 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 16114 12724 16120 12776
rect 16172 12724 16178 12776
rect 16485 12767 16543 12773
rect 16485 12733 16497 12767
rect 16531 12764 16543 12767
rect 16574 12764 16580 12776
rect 16531 12736 16580 12764
rect 16531 12733 16543 12736
rect 16485 12727 16543 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 16684 12773 16712 12804
rect 16758 12792 16764 12844
rect 16816 12832 16822 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16816 12804 16957 12832
rect 16816 12792 16822 12804
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 16945 12795 17003 12801
rect 17402 12792 17408 12844
rect 17460 12792 17466 12844
rect 17604 12832 17632 12872
rect 18325 12869 18337 12872
rect 18371 12869 18383 12903
rect 18325 12863 18383 12869
rect 18414 12832 18420 12844
rect 17512 12804 17632 12832
rect 17788 12804 18420 12832
rect 16669 12767 16727 12773
rect 16669 12733 16681 12767
rect 16715 12733 16727 12767
rect 16669 12727 16727 12733
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12733 16911 12767
rect 16853 12727 16911 12733
rect 14829 12699 14887 12705
rect 14829 12696 14841 12699
rect 14768 12668 14841 12696
rect 14829 12665 14841 12668
rect 14875 12665 14887 12699
rect 14829 12659 14887 12665
rect 14921 12699 14979 12705
rect 14921 12665 14933 12699
rect 14967 12696 14979 12699
rect 16022 12696 16028 12708
rect 14967 12668 16028 12696
rect 14967 12665 14979 12668
rect 14921 12659 14979 12665
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 16132 12696 16160 12724
rect 16868 12696 16896 12727
rect 17034 12724 17040 12776
rect 17092 12724 17098 12776
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12764 17187 12767
rect 17512 12764 17540 12804
rect 17788 12773 17816 12804
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 17175 12736 17540 12764
rect 17773 12767 17831 12773
rect 17175 12733 17187 12736
rect 17129 12727 17187 12733
rect 17773 12733 17785 12767
rect 17819 12733 17831 12767
rect 17773 12727 17831 12733
rect 16132 12668 16896 12696
rect 6043 12600 6408 12628
rect 6733 12631 6791 12637
rect 6043 12597 6055 12600
rect 5997 12591 6055 12597
rect 6733 12597 6745 12631
rect 6779 12597 6791 12631
rect 6733 12591 6791 12597
rect 6914 12588 6920 12640
rect 6972 12588 6978 12640
rect 10689 12631 10747 12637
rect 10689 12597 10701 12631
rect 10735 12628 10747 12631
rect 11974 12628 11980 12640
rect 10735 12600 11980 12628
rect 10735 12597 10747 12600
rect 10689 12591 10747 12597
rect 11974 12588 11980 12600
rect 12032 12588 12038 12640
rect 14734 12588 14740 12640
rect 14792 12628 14798 12640
rect 15105 12631 15163 12637
rect 15105 12628 15117 12631
rect 14792 12600 15117 12628
rect 14792 12588 14798 12600
rect 15105 12597 15117 12600
rect 15151 12597 15163 12631
rect 15105 12591 15163 12597
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15565 12631 15623 12637
rect 15565 12628 15577 12631
rect 15252 12600 15577 12628
rect 15252 12588 15258 12600
rect 15565 12597 15577 12600
rect 15611 12597 15623 12631
rect 15565 12591 15623 12597
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 17144 12628 17172 12727
rect 17586 12637 17592 12640
rect 15712 12600 17172 12628
rect 17570 12631 17592 12637
rect 15712 12588 15718 12600
rect 17570 12597 17582 12631
rect 17570 12591 17592 12597
rect 17586 12588 17592 12591
rect 17644 12588 17650 12640
rect 17678 12588 17684 12640
rect 17736 12588 17742 12640
rect 1104 12538 18860 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 18860 12538
rect 1104 12464 18860 12486
rect 1578 12384 1584 12436
rect 1636 12384 1642 12436
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12424 3663 12427
rect 3786 12424 3792 12436
rect 3651 12396 3792 12424
rect 3651 12393 3663 12396
rect 3605 12387 3663 12393
rect 3786 12384 3792 12396
rect 3844 12384 3850 12436
rect 5077 12427 5135 12433
rect 5077 12393 5089 12427
rect 5123 12424 5135 12427
rect 5350 12424 5356 12436
rect 5123 12396 5356 12424
rect 5123 12393 5135 12396
rect 5077 12387 5135 12393
rect 2498 12316 2504 12368
rect 2556 12356 2562 12368
rect 2593 12359 2651 12365
rect 2593 12356 2605 12359
rect 2556 12328 2605 12356
rect 2556 12316 2562 12328
rect 2593 12325 2605 12328
rect 2639 12325 2651 12359
rect 2593 12319 2651 12325
rect 3418 12316 3424 12368
rect 3476 12356 3482 12368
rect 3476 12328 4292 12356
rect 3476 12316 3482 12328
rect 1670 12248 1676 12300
rect 1728 12288 1734 12300
rect 4154 12288 4160 12300
rect 1728 12260 3372 12288
rect 1728 12248 1734 12260
rect 842 12180 848 12232
rect 900 12220 906 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 900 12192 1409 12220
rect 900 12180 906 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2222 12220 2228 12232
rect 2179 12192 2228 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2222 12180 2228 12192
rect 2280 12180 2286 12232
rect 2424 12229 2452 12260
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12189 2467 12223
rect 2409 12183 2467 12189
rect 2590 12180 2596 12232
rect 2648 12214 2654 12232
rect 2685 12223 2743 12229
rect 2685 12214 2697 12223
rect 2648 12189 2697 12214
rect 2731 12189 2743 12223
rect 2648 12186 2743 12189
rect 2648 12180 2654 12186
rect 2685 12183 2743 12186
rect 2869 12223 2927 12229
rect 2869 12189 2881 12223
rect 2915 12189 2927 12223
rect 2869 12183 2927 12189
rect 2498 12112 2504 12164
rect 2556 12152 2562 12164
rect 2884 12152 2912 12183
rect 2556 12124 2912 12152
rect 3237 12155 3295 12161
rect 2556 12112 2562 12124
rect 3237 12121 3249 12155
rect 3283 12121 3295 12155
rect 3344 12152 3372 12260
rect 3528 12260 4160 12288
rect 3418 12180 3424 12232
rect 3476 12180 3482 12232
rect 3528 12152 3556 12260
rect 4154 12248 4160 12260
rect 4212 12248 4218 12300
rect 4264 12297 4292 12328
rect 4249 12291 4307 12297
rect 4249 12257 4261 12291
rect 4295 12288 4307 12291
rect 4295 12260 4936 12288
rect 4295 12257 4307 12260
rect 4249 12251 4307 12257
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 3344 12124 3556 12152
rect 3896 12152 3924 12183
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 4028 12192 4077 12220
rect 4028 12180 4034 12192
rect 4065 12189 4077 12192
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 4430 12180 4436 12232
rect 4488 12220 4494 12232
rect 4706 12220 4712 12232
rect 4488 12192 4712 12220
rect 4488 12180 4494 12192
rect 4706 12180 4712 12192
rect 4764 12180 4770 12232
rect 4908 12229 4936 12260
rect 4893 12223 4951 12229
rect 4893 12189 4905 12223
rect 4939 12220 4951 12223
rect 4982 12220 4988 12232
rect 4939 12192 4988 12220
rect 4939 12189 4951 12192
rect 4893 12183 4951 12189
rect 4982 12180 4988 12192
rect 5040 12180 5046 12232
rect 5184 12229 5212 12396
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 7248 12396 8217 12424
rect 7248 12384 7254 12396
rect 8205 12393 8217 12396
rect 8251 12393 8263 12427
rect 8205 12387 8263 12393
rect 10505 12427 10563 12433
rect 10505 12393 10517 12427
rect 10551 12424 10563 12427
rect 10686 12424 10692 12436
rect 10551 12396 10692 12424
rect 10551 12393 10563 12396
rect 10505 12387 10563 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 14458 12384 14464 12436
rect 14516 12384 14522 12436
rect 15930 12424 15936 12436
rect 14752 12396 15936 12424
rect 5350 12248 5356 12300
rect 5408 12288 5414 12300
rect 5445 12291 5503 12297
rect 5445 12288 5457 12291
rect 5408 12260 5457 12288
rect 5408 12248 5414 12260
rect 5445 12257 5457 12260
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 7926 12248 7932 12300
rect 7984 12288 7990 12300
rect 7984 12260 8524 12288
rect 7984 12248 7990 12260
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 5261 12223 5319 12229
rect 5261 12189 5273 12223
rect 5307 12189 5319 12223
rect 5261 12183 5319 12189
rect 4617 12155 4675 12161
rect 3896 12124 4568 12152
rect 3237 12115 3295 12121
rect 2225 12087 2283 12093
rect 2225 12053 2237 12087
rect 2271 12084 2283 12087
rect 2958 12084 2964 12096
rect 2271 12056 2964 12084
rect 2271 12053 2283 12056
rect 2225 12047 2283 12053
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 3053 12087 3111 12093
rect 3053 12053 3065 12087
rect 3099 12084 3111 12087
rect 3252 12084 3280 12115
rect 3970 12084 3976 12096
rect 3099 12056 3976 12084
rect 3099 12053 3111 12056
rect 3053 12047 3111 12053
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4540 12084 4568 12124
rect 4617 12121 4629 12155
rect 4663 12152 4675 12155
rect 5276 12152 5304 12183
rect 6454 12180 6460 12232
rect 6512 12180 6518 12232
rect 8496 12229 8524 12260
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10689 12291 10747 12297
rect 10689 12288 10701 12291
rect 9732 12260 10701 12288
rect 9732 12248 9738 12260
rect 10689 12257 10701 12260
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 14642 12248 14648 12300
rect 14700 12248 14706 12300
rect 14752 12297 14780 12396
rect 15930 12384 15936 12396
rect 15988 12424 15994 12436
rect 16114 12424 16120 12436
rect 15988 12396 16120 12424
rect 15988 12384 15994 12396
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17092 12396 17509 12424
rect 17092 12384 17098 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 17497 12387 17555 12393
rect 15102 12316 15108 12368
rect 15160 12316 15166 12368
rect 17052 12356 17080 12384
rect 15488 12328 17080 12356
rect 18325 12359 18383 12365
rect 14737 12291 14795 12297
rect 14737 12257 14749 12291
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12288 14979 12291
rect 15194 12288 15200 12300
rect 14967 12260 15200 12288
rect 14967 12257 14979 12260
rect 14921 12251 14979 12257
rect 15194 12248 15200 12260
rect 15252 12248 15258 12300
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 4663 12124 5304 12152
rect 6733 12155 6791 12161
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 6733 12121 6745 12155
rect 6779 12152 6791 12155
rect 8389 12155 8447 12161
rect 8389 12152 8401 12155
rect 6779 12124 6960 12152
rect 7958 12124 8401 12152
rect 6779 12121 6791 12124
rect 6733 12115 6791 12121
rect 6932 12096 6960 12124
rect 8389 12121 8401 12124
rect 8435 12121 8447 12155
rect 8496 12152 8524 12183
rect 9858 12180 9864 12232
rect 9916 12220 9922 12232
rect 10045 12223 10103 12229
rect 10045 12220 10057 12223
rect 9916 12192 10057 12220
rect 9916 12180 9922 12192
rect 10045 12189 10057 12192
rect 10091 12189 10103 12223
rect 10045 12183 10103 12189
rect 10134 12180 10140 12232
rect 10192 12180 10198 12232
rect 10321 12223 10379 12229
rect 10321 12189 10333 12223
rect 10367 12220 10379 12223
rect 10502 12220 10508 12232
rect 10367 12192 10508 12220
rect 10367 12189 10379 12192
rect 10321 12183 10379 12189
rect 10502 12180 10508 12192
rect 10560 12180 10566 12232
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12220 11299 12223
rect 11330 12220 11336 12232
rect 11287 12192 11336 12220
rect 11287 12189 11299 12192
rect 11241 12183 11299 12189
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 11808 12152 11836 12183
rect 8496 12124 11836 12152
rect 8389 12115 8447 12121
rect 5258 12084 5264 12096
rect 4540 12056 5264 12084
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 5442 12044 5448 12096
rect 5500 12044 5506 12096
rect 6914 12044 6920 12096
rect 6972 12044 6978 12096
rect 11882 12044 11888 12096
rect 11940 12044 11946 12096
rect 14844 12084 14872 12183
rect 15010 12180 15016 12232
rect 15068 12220 15074 12232
rect 15488 12229 15516 12328
rect 18325 12325 18337 12359
rect 18371 12325 18383 12359
rect 18325 12319 18383 12325
rect 15565 12291 15623 12297
rect 15565 12257 15577 12291
rect 15611 12288 15623 12291
rect 15654 12288 15660 12300
rect 15611 12260 15660 12288
rect 15611 12257 15623 12260
rect 15565 12251 15623 12257
rect 15654 12248 15660 12260
rect 15712 12248 15718 12300
rect 15473 12223 15531 12229
rect 15473 12220 15485 12223
rect 15068 12192 15485 12220
rect 15068 12180 15074 12192
rect 15473 12189 15485 12192
rect 15519 12189 15531 12223
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 15473 12183 15531 12189
rect 15672 12192 15761 12220
rect 15672 12084 15700 12192
rect 15749 12189 15761 12192
rect 15795 12220 15807 12223
rect 15795 12192 15884 12220
rect 15795 12189 15807 12192
rect 15749 12183 15807 12189
rect 15856 12152 15884 12192
rect 15930 12180 15936 12232
rect 15988 12180 15994 12232
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 17402 12220 17408 12232
rect 16080 12192 17408 12220
rect 16080 12180 16086 12192
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12220 17647 12223
rect 17678 12220 17684 12232
rect 17635 12192 17684 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 17678 12180 17684 12192
rect 17736 12220 17742 12232
rect 18340 12220 18368 12319
rect 17736 12192 18368 12220
rect 17736 12180 17742 12192
rect 18506 12180 18512 12232
rect 18564 12180 18570 12232
rect 16758 12152 16764 12164
rect 15856 12124 16764 12152
rect 16758 12112 16764 12124
rect 16816 12112 16822 12164
rect 14844 12056 15700 12084
rect 15746 12044 15752 12096
rect 15804 12044 15810 12096
rect 1104 11994 18860 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 18860 11994
rect 1104 11920 18860 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 2038 11880 2044 11892
rect 1627 11852 2044 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 2038 11840 2044 11852
rect 2096 11840 2102 11892
rect 2682 11840 2688 11892
rect 2740 11880 2746 11892
rect 4430 11880 4436 11892
rect 2740 11852 4436 11880
rect 2740 11840 2746 11852
rect 4430 11840 4436 11852
rect 4488 11840 4494 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 7561 11883 7619 11889
rect 7561 11880 7573 11883
rect 5500 11852 7573 11880
rect 5500 11840 5506 11852
rect 7561 11849 7573 11852
rect 7607 11849 7619 11883
rect 12526 11880 12532 11892
rect 7561 11843 7619 11849
rect 9876 11852 12532 11880
rect 7926 11812 7932 11824
rect 2746 11784 7932 11812
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 900 11716 1409 11744
rect 900 11704 906 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2225 11747 2283 11753
rect 2225 11713 2237 11747
rect 2271 11744 2283 11747
rect 2746 11744 2774 11784
rect 7926 11772 7932 11784
rect 7984 11772 7990 11824
rect 8018 11772 8024 11824
rect 8076 11772 8082 11824
rect 9582 11772 9588 11824
rect 9640 11772 9646 11824
rect 9876 11756 9904 11852
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 11790 11812 11796 11824
rect 10827 11784 11796 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 11940 11784 12282 11812
rect 13372 11784 14320 11812
rect 11940 11772 11946 11784
rect 2271 11716 2774 11744
rect 3973 11747 4031 11753
rect 2271 11713 2283 11716
rect 2225 11707 2283 11713
rect 3973 11713 3985 11747
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 1578 11636 1584 11688
rect 1636 11676 1642 11688
rect 3988 11676 4016 11707
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 4120 11716 4165 11744
rect 4120 11704 4126 11716
rect 9858 11704 9864 11756
rect 9916 11704 9922 11756
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11744 10103 11747
rect 10134 11744 10140 11756
rect 10091 11716 10140 11744
rect 10091 11713 10103 11716
rect 10045 11707 10103 11713
rect 10134 11704 10140 11716
rect 10192 11704 10198 11756
rect 10870 11704 10876 11756
rect 10928 11744 10934 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10928 11716 11529 11744
rect 10928 11704 10934 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 4614 11676 4620 11688
rect 1636 11648 4620 11676
rect 1636 11636 1642 11648
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10413 11679 10471 11685
rect 10413 11676 10425 11679
rect 10008 11648 10425 11676
rect 10008 11636 10014 11648
rect 10413 11645 10425 11648
rect 10459 11676 10471 11679
rect 10778 11676 10784 11688
rect 10459 11648 10784 11676
rect 10459 11645 10471 11648
rect 10413 11639 10471 11645
rect 10778 11636 10784 11648
rect 10836 11636 10842 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 10980 11648 11805 11676
rect 7377 11611 7435 11617
rect 7377 11577 7389 11611
rect 7423 11608 7435 11611
rect 7929 11611 7987 11617
rect 7423 11580 7880 11608
rect 7423 11577 7435 11580
rect 7377 11571 7435 11577
rect 2130 11500 2136 11552
rect 2188 11500 2194 11552
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 5534 11540 5540 11552
rect 4203 11512 5540 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 5534 11500 5540 11512
rect 5592 11540 5598 11552
rect 7561 11543 7619 11549
rect 7561 11540 7573 11543
rect 5592 11512 7573 11540
rect 5592 11500 5598 11512
rect 7561 11509 7573 11512
rect 7607 11509 7619 11543
rect 7852 11540 7880 11580
rect 7929 11577 7941 11611
rect 7975 11608 7987 11611
rect 9122 11608 9128 11620
rect 7975 11580 9128 11608
rect 7975 11577 7987 11580
rect 7929 11571 7987 11577
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 10980 11617 11008 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 11793 11639 11851 11645
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13372 11685 13400 11784
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13587 11716 13829 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 13357 11679 13415 11685
rect 13357 11676 13369 11679
rect 13320 11648 13369 11676
rect 13320 11636 13326 11648
rect 13357 11645 13369 11648
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 10965 11611 11023 11617
rect 10965 11577 10977 11611
rect 11011 11577 11023 11611
rect 10965 11571 11023 11577
rect 13648 11608 13676 11716
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 13998 11704 14004 11756
rect 14056 11704 14062 11756
rect 14090 11704 14096 11756
rect 14148 11704 14154 11756
rect 14292 11753 14320 11784
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 13725 11679 13783 11685
rect 13725 11645 13737 11679
rect 13771 11676 13783 11679
rect 14016 11676 14044 11704
rect 13771 11648 14044 11676
rect 15580 11676 15608 11707
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16850 11744 16856 11756
rect 15887 11716 16856 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 16942 11676 16948 11688
rect 15580 11648 16948 11676
rect 13771 11645 13783 11648
rect 13725 11639 13783 11645
rect 15580 11608 15608 11648
rect 16942 11636 16948 11648
rect 17000 11636 17006 11688
rect 13648 11580 15608 11608
rect 8938 11540 8944 11552
rect 7852 11512 8944 11540
rect 7561 11503 7619 11509
rect 8938 11500 8944 11512
rect 8996 11500 9002 11552
rect 9306 11500 9312 11552
rect 9364 11540 9370 11552
rect 9953 11543 10011 11549
rect 9953 11540 9965 11543
rect 9364 11512 9965 11540
rect 9364 11500 9370 11512
rect 9953 11509 9965 11512
rect 9999 11509 10011 11543
rect 9953 11503 10011 11509
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 10781 11543 10839 11549
rect 10781 11540 10793 11543
rect 10284 11512 10793 11540
rect 10284 11500 10290 11512
rect 10781 11509 10793 11512
rect 10827 11509 10839 11543
rect 10781 11503 10839 11509
rect 13265 11543 13323 11549
rect 13265 11509 13277 11543
rect 13311 11540 13323 11543
rect 13538 11540 13544 11552
rect 13311 11512 13544 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 13538 11500 13544 11512
rect 13596 11540 13602 11552
rect 13648 11540 13676 11580
rect 13596 11512 13676 11540
rect 13596 11500 13602 11512
rect 13814 11500 13820 11552
rect 13872 11500 13878 11552
rect 13906 11500 13912 11552
rect 13964 11540 13970 11552
rect 14093 11543 14151 11549
rect 14093 11540 14105 11543
rect 13964 11512 14105 11540
rect 13964 11500 13970 11512
rect 14093 11509 14105 11512
rect 14139 11509 14151 11543
rect 14093 11503 14151 11509
rect 15378 11500 15384 11552
rect 15436 11500 15442 11552
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 16758 11540 16764 11552
rect 16080 11512 16764 11540
rect 16080 11500 16086 11512
rect 16758 11500 16764 11512
rect 16816 11500 16822 11552
rect 1104 11450 18860 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 18860 11450
rect 1104 11376 18860 11398
rect 1394 11296 1400 11348
rect 1452 11296 1458 11348
rect 4617 11339 4675 11345
rect 4617 11305 4629 11339
rect 4663 11336 4675 11339
rect 5350 11336 5356 11348
rect 4663 11308 5356 11336
rect 4663 11305 4675 11308
rect 4617 11299 4675 11305
rect 5350 11296 5356 11308
rect 5408 11296 5414 11348
rect 5534 11296 5540 11348
rect 5592 11296 5598 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 5920 11308 8953 11336
rect 5920 11268 5948 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 10778 11296 10784 11348
rect 10836 11296 10842 11348
rect 11790 11296 11796 11348
rect 11848 11296 11854 11348
rect 13909 11339 13967 11345
rect 13909 11305 13921 11339
rect 13955 11336 13967 11339
rect 14090 11336 14096 11348
rect 13955 11308 14096 11336
rect 13955 11305 13967 11308
rect 13909 11299 13967 11305
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 15746 11296 15752 11348
rect 15804 11336 15810 11348
rect 16761 11339 16819 11345
rect 16761 11336 16773 11339
rect 15804 11308 16773 11336
rect 15804 11296 15810 11308
rect 16761 11305 16773 11308
rect 16807 11305 16819 11339
rect 16761 11299 16819 11305
rect 3068 11240 5948 11268
rect 2869 11203 2927 11209
rect 2869 11169 2881 11203
rect 2915 11200 2927 11203
rect 3068 11200 3096 11240
rect 8570 11228 8576 11280
rect 8628 11268 8634 11280
rect 9217 11271 9275 11277
rect 9217 11268 9229 11271
rect 8628 11240 9229 11268
rect 8628 11228 8634 11240
rect 9217 11237 9229 11240
rect 9263 11237 9275 11271
rect 12894 11268 12900 11280
rect 9217 11231 9275 11237
rect 9784 11240 12900 11268
rect 2915 11172 3096 11200
rect 3145 11203 3203 11209
rect 2915 11169 2927 11172
rect 2869 11163 2927 11169
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 5813 11203 5871 11209
rect 5813 11200 5825 11203
rect 3191 11172 5825 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 5813 11169 5825 11172
rect 5859 11200 5871 11203
rect 6454 11200 6460 11212
rect 5859 11172 6460 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6546 11160 6552 11212
rect 6604 11200 6610 11212
rect 7561 11203 7619 11209
rect 7561 11200 7573 11203
rect 6604 11172 7573 11200
rect 6604 11160 6610 11172
rect 7561 11169 7573 11172
rect 7607 11169 7619 11203
rect 7561 11163 7619 11169
rect 9306 11160 9312 11212
rect 9364 11160 9370 11212
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9447 11172 9689 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 3418 11092 3424 11144
rect 3476 11132 3482 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3476 11104 3801 11132
rect 3476 11092 3482 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4246 11132 4252 11144
rect 4203 11104 4252 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4246 11092 4252 11104
rect 4304 11092 4310 11144
rect 4430 11092 4436 11144
rect 4488 11092 4494 11144
rect 4614 11141 4620 11144
rect 4587 11135 4620 11141
rect 4587 11101 4599 11135
rect 4587 11095 4620 11101
rect 4614 11092 4620 11095
rect 4672 11092 4678 11144
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5350 11132 5356 11144
rect 5215 11104 5356 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 7926 11092 7932 11144
rect 7984 11092 7990 11144
rect 9122 11092 9128 11144
rect 9180 11092 9186 11144
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 9784 11132 9812 11240
rect 12894 11228 12900 11240
rect 12952 11228 12958 11280
rect 16298 11268 16304 11280
rect 16224 11240 16304 11268
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11200 10195 11203
rect 13906 11200 13912 11212
rect 10183 11172 13912 11200
rect 10183 11169 10195 11172
rect 10137 11163 10195 11169
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 16224 11209 16252 11240
rect 16298 11228 16304 11240
rect 16356 11228 16362 11280
rect 16577 11271 16635 11277
rect 16577 11268 16589 11271
rect 16408 11240 16589 11268
rect 16408 11209 16436 11240
rect 16577 11237 16589 11240
rect 16623 11237 16635 11271
rect 16577 11231 16635 11237
rect 16209 11203 16267 11209
rect 16209 11169 16221 11203
rect 16255 11169 16267 11203
rect 16209 11163 16267 11169
rect 16393 11203 16451 11209
rect 16393 11169 16405 11203
rect 16439 11169 16451 11203
rect 16393 11163 16451 11169
rect 9631 11104 9812 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 10042 11092 10048 11144
rect 10100 11092 10106 11144
rect 10413 11135 10471 11141
rect 10413 11101 10425 11135
rect 10459 11101 10471 11135
rect 10413 11095 10471 11101
rect 2130 11024 2136 11076
rect 2188 11024 2194 11076
rect 4062 11024 4068 11076
rect 4120 11064 4126 11076
rect 4448 11064 4476 11092
rect 4120 11036 4476 11064
rect 5537 11067 5595 11073
rect 4120 11024 4126 11036
rect 5537 11033 5549 11067
rect 5583 11064 5595 11067
rect 5626 11064 5632 11076
rect 5583 11036 5632 11064
rect 5583 11033 5595 11036
rect 5537 11027 5595 11033
rect 5626 11024 5632 11036
rect 5684 11024 5690 11076
rect 6089 11067 6147 11073
rect 6089 11064 6101 11067
rect 5736 11036 6101 11064
rect 4154 10956 4160 11008
rect 4212 10996 4218 11008
rect 5736 11005 5764 11036
rect 6089 11033 6101 11036
rect 6135 11033 6147 11067
rect 7837 11067 7895 11073
rect 7837 11064 7849 11067
rect 7314 11036 7849 11064
rect 6089 11027 6147 11033
rect 7837 11033 7849 11036
rect 7883 11033 7895 11067
rect 7837 11027 7895 11033
rect 8662 11024 8668 11076
rect 8720 11064 8726 11076
rect 9398 11064 9404 11076
rect 8720 11036 9404 11064
rect 8720 11024 8726 11036
rect 9398 11024 9404 11036
rect 9456 11064 9462 11076
rect 10428 11064 10456 11095
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 11020 11104 11069 11132
rect 11020 11092 11026 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 11333 11135 11391 11141
rect 11333 11101 11345 11135
rect 11379 11132 11391 11135
rect 11379 11104 11652 11132
rect 11379 11101 11391 11104
rect 11333 11095 11391 11101
rect 11238 11064 11244 11076
rect 9456 11036 10456 11064
rect 10612 11036 11244 11064
rect 9456 11024 9462 11036
rect 10612 11005 10640 11036
rect 11238 11024 11244 11036
rect 11296 11024 11302 11076
rect 11422 11024 11428 11076
rect 11480 11024 11486 11076
rect 11624 11073 11652 11104
rect 13170 11092 13176 11144
rect 13228 11092 13234 11144
rect 13354 11092 13360 11144
rect 13412 11092 13418 11144
rect 13446 11092 13452 11144
rect 13504 11092 13510 11144
rect 13538 11092 13544 11144
rect 13596 11092 13602 11144
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 13998 11132 14004 11144
rect 13771 11104 14004 11132
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 13998 11092 14004 11104
rect 14056 11092 14062 11144
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 15838 11132 15844 11144
rect 15344 11104 15844 11132
rect 15344 11092 15350 11104
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 16301 11135 16359 11141
rect 16301 11101 16313 11135
rect 16347 11132 16359 11135
rect 17865 11135 17923 11141
rect 16347 11104 16528 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 11609 11067 11667 11073
rect 11609 11033 11621 11067
rect 11655 11064 11667 11067
rect 13556 11064 13584 11092
rect 16132 11064 16160 11095
rect 16390 11064 16396 11076
rect 11655 11036 13584 11064
rect 15856 11036 16068 11064
rect 16132 11036 16396 11064
rect 11655 11033 11667 11036
rect 11609 11027 11667 11033
rect 4341 10999 4399 11005
rect 4341 10996 4353 10999
rect 4212 10968 4353 10996
rect 4212 10956 4218 10968
rect 4341 10965 4353 10968
rect 4387 10965 4399 10999
rect 4341 10959 4399 10965
rect 5721 10999 5779 11005
rect 5721 10965 5733 10999
rect 5767 10965 5779 10999
rect 5721 10959 5779 10965
rect 10597 10999 10655 11005
rect 10597 10965 10609 10999
rect 10643 10965 10655 10999
rect 10597 10959 10655 10965
rect 10686 10956 10692 11008
rect 10744 10996 10750 11008
rect 10965 10999 11023 11005
rect 10965 10996 10977 10999
rect 10744 10968 10977 10996
rect 10744 10956 10750 10968
rect 10965 10965 10977 10968
rect 11011 10965 11023 10999
rect 10965 10959 11023 10965
rect 11146 10956 11152 11008
rect 11204 10996 11210 11008
rect 12342 10996 12348 11008
rect 11204 10968 12348 10996
rect 11204 10956 11210 10968
rect 12342 10956 12348 10968
rect 12400 10996 12406 11008
rect 15856 10996 15884 11036
rect 12400 10968 15884 10996
rect 12400 10956 12406 10968
rect 15930 10956 15936 11008
rect 15988 10956 15994 11008
rect 16040 10996 16068 11036
rect 16390 11024 16396 11036
rect 16448 11024 16454 11076
rect 16114 10996 16120 11008
rect 16040 10968 16120 10996
rect 16114 10956 16120 10968
rect 16172 10996 16178 11008
rect 16500 10996 16528 11104
rect 17865 11101 17877 11135
rect 17911 11132 17923 11135
rect 17911 11104 18092 11132
rect 17911 11101 17923 11104
rect 17865 11095 17923 11101
rect 16745 11067 16803 11073
rect 16745 11033 16757 11067
rect 16791 11064 16803 11067
rect 16850 11064 16856 11076
rect 16791 11036 16856 11064
rect 16791 11033 16803 11036
rect 16745 11027 16803 11033
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 16942 11024 16948 11076
rect 17000 11024 17006 11076
rect 16172 10968 16528 10996
rect 16172 10956 16178 10968
rect 17218 10956 17224 11008
rect 17276 10996 17282 11008
rect 17773 10999 17831 11005
rect 17773 10996 17785 10999
rect 17276 10968 17785 10996
rect 17276 10956 17282 10968
rect 17773 10965 17785 10968
rect 17819 10965 17831 10999
rect 17773 10959 17831 10965
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18064 11005 18092 11104
rect 18230 11092 18236 11144
rect 18288 11092 18294 11144
rect 18506 11092 18512 11144
rect 18564 11092 18570 11144
rect 18049 10999 18107 11005
rect 18049 10996 18061 10999
rect 18012 10968 18061 10996
rect 18012 10956 18018 10968
rect 18049 10965 18061 10968
rect 18095 10965 18107 10999
rect 18049 10959 18107 10965
rect 18322 10956 18328 11008
rect 18380 10956 18386 11008
rect 1104 10906 18860 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 18860 10906
rect 1104 10832 18860 10854
rect 1578 10752 1584 10804
rect 1636 10752 1642 10804
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 4246 10792 4252 10804
rect 2823 10764 4252 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 4246 10752 4252 10764
rect 4304 10752 4310 10804
rect 5534 10752 5540 10804
rect 5592 10752 5598 10804
rect 9217 10795 9275 10801
rect 9217 10761 9229 10795
rect 9263 10792 9275 10795
rect 10042 10792 10048 10804
rect 9263 10764 10048 10792
rect 9263 10761 9275 10764
rect 9217 10755 9275 10761
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 11149 10795 11207 10801
rect 11149 10792 11161 10795
rect 10336 10764 11161 10792
rect 4706 10724 4712 10736
rect 3988 10696 4712 10724
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 900 10628 1409 10656
rect 900 10616 906 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 2409 10659 2467 10665
rect 2409 10625 2421 10659
rect 2455 10656 2467 10659
rect 2682 10656 2688 10668
rect 2455 10628 2688 10656
rect 2455 10625 2467 10628
rect 2409 10619 2467 10625
rect 2682 10616 2688 10628
rect 2740 10616 2746 10668
rect 3988 10665 4016 10696
rect 4706 10684 4712 10696
rect 4764 10684 4770 10736
rect 5442 10724 5448 10736
rect 5276 10696 5448 10724
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 4433 10659 4491 10665
rect 4433 10625 4445 10659
rect 4479 10656 4491 10659
rect 4798 10656 4804 10668
rect 4479 10628 4804 10656
rect 4479 10625 4491 10628
rect 4433 10619 4491 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 5276 10665 5304 10696
rect 5442 10684 5448 10696
rect 5500 10724 5506 10736
rect 5902 10724 5908 10736
rect 5500 10696 5908 10724
rect 5500 10684 5506 10696
rect 5902 10684 5908 10696
rect 5960 10684 5966 10736
rect 6546 10724 6552 10736
rect 6012 10696 6552 10724
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10625 5319 10659
rect 5261 10619 5319 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 6012 10656 6040 10696
rect 6546 10684 6552 10696
rect 6604 10684 6610 10736
rect 9674 10684 9680 10736
rect 9732 10684 9738 10736
rect 5767 10628 6040 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2590 10588 2596 10600
rect 2547 10560 2596 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2590 10548 2596 10560
rect 2648 10548 2654 10600
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 4522 10588 4528 10600
rect 3936 10560 4528 10588
rect 3936 10548 3942 10560
rect 4522 10548 4528 10560
rect 4580 10588 4586 10600
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 4580 10560 5089 10588
rect 4580 10548 4586 10560
rect 5077 10557 5089 10560
rect 5123 10588 5135 10591
rect 5736 10588 5764 10619
rect 7742 10616 7748 10668
rect 7800 10616 7806 10668
rect 8757 10659 8815 10665
rect 8757 10625 8769 10659
rect 8803 10625 8815 10659
rect 8757 10619 8815 10625
rect 5123 10560 5764 10588
rect 6365 10591 6423 10597
rect 5123 10557 5135 10560
rect 5077 10551 5135 10557
rect 6365 10557 6377 10591
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 4617 10455 4675 10461
rect 4617 10421 4629 10455
rect 4663 10452 4675 10455
rect 5258 10452 5264 10464
rect 4663 10424 5264 10452
rect 4663 10421 4675 10424
rect 4617 10415 4675 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 5408 10424 5457 10452
rect 5408 10412 5414 10424
rect 5445 10421 5457 10424
rect 5491 10421 5503 10455
rect 6380 10452 6408 10551
rect 6638 10548 6644 10600
rect 6696 10548 6702 10600
rect 8772 10588 8800 10619
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 10045 10659 10103 10665
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10336 10656 10364 10764
rect 11149 10761 11161 10764
rect 11195 10792 11207 10795
rect 11422 10792 11428 10804
rect 11195 10764 11428 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 11422 10752 11428 10764
rect 11480 10752 11486 10804
rect 12989 10795 13047 10801
rect 12989 10761 13001 10795
rect 13035 10792 13047 10795
rect 13170 10792 13176 10804
rect 13035 10764 13176 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 13446 10752 13452 10804
rect 13504 10792 13510 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 13504 10764 13737 10792
rect 13504 10752 13510 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 13725 10755 13783 10761
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 14700 10764 16620 10792
rect 14700 10752 14706 10764
rect 10781 10727 10839 10733
rect 10781 10724 10793 10727
rect 10428 10696 10793 10724
rect 10428 10665 10456 10696
rect 10781 10693 10793 10696
rect 10827 10693 10839 10727
rect 10781 10687 10839 10693
rect 10091 10628 10364 10656
rect 10413 10659 10471 10665
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10413 10625 10425 10659
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 10597 10659 10655 10665
rect 10597 10625 10609 10659
rect 10643 10625 10655 10659
rect 10597 10619 10655 10625
rect 10134 10588 10140 10600
rect 8772 10560 10140 10588
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 10612 10588 10640 10619
rect 10686 10616 10692 10668
rect 10744 10616 10750 10668
rect 10796 10656 10824 10687
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 10981 10727 11039 10733
rect 10981 10724 10993 10727
rect 10928 10696 10993 10724
rect 10928 10684 10934 10696
rect 10981 10693 10993 10696
rect 11027 10693 11039 10727
rect 12805 10727 12863 10733
rect 12805 10724 12817 10727
rect 10981 10687 11039 10693
rect 12176 10696 12817 10724
rect 11146 10656 11152 10668
rect 10796 10628 11152 10656
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 12176 10665 12204 10696
rect 12805 10693 12817 10696
rect 12851 10724 12863 10727
rect 15010 10724 15016 10736
rect 12851 10696 15016 10724
rect 12851 10693 12863 10696
rect 12805 10687 12863 10693
rect 15010 10684 15016 10696
rect 15068 10684 15074 10736
rect 15194 10724 15200 10736
rect 15120 10696 15200 10724
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10625 12219 10659
rect 12342 10656 12348 10668
rect 12303 10628 12348 10656
rect 12161 10619 12219 10625
rect 12342 10616 12348 10628
rect 12400 10656 12406 10668
rect 12621 10659 12679 10665
rect 12621 10656 12633 10659
rect 12400 10628 12633 10656
rect 12400 10616 12406 10628
rect 12621 10625 12633 10628
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 13170 10616 13176 10668
rect 13228 10656 13234 10668
rect 13633 10659 13691 10665
rect 13633 10656 13645 10659
rect 13228 10628 13645 10656
rect 13228 10616 13234 10628
rect 13633 10625 13645 10628
rect 13679 10625 13691 10659
rect 13633 10619 13691 10625
rect 13909 10659 13967 10665
rect 13909 10625 13921 10659
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 13357 10591 13415 10597
rect 10612 10560 11008 10588
rect 8846 10480 8852 10532
rect 8904 10480 8910 10532
rect 10980 10464 11008 10560
rect 13357 10557 13369 10591
rect 13403 10588 13415 10591
rect 13814 10588 13820 10600
rect 13403 10560 13820 10588
rect 13403 10557 13415 10560
rect 13357 10551 13415 10557
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 12529 10523 12587 10529
rect 12529 10489 12541 10523
rect 12575 10520 12587 10523
rect 12575 10492 13400 10520
rect 12575 10489 12587 10492
rect 12529 10483 12587 10489
rect 13372 10464 13400 10492
rect 7098 10452 7104 10464
rect 6380 10424 7104 10452
rect 5445 10415 5503 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 9490 10412 9496 10464
rect 9548 10412 9554 10464
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 10229 10455 10287 10461
rect 10229 10452 10241 10455
rect 9723 10424 10241 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 10229 10421 10241 10424
rect 10275 10421 10287 10455
rect 10229 10415 10287 10421
rect 10962 10412 10968 10464
rect 11020 10412 11026 10464
rect 13078 10412 13084 10464
rect 13136 10412 13142 10464
rect 13354 10412 13360 10464
rect 13412 10412 13418 10464
rect 13541 10455 13599 10461
rect 13541 10421 13553 10455
rect 13587 10452 13599 10455
rect 13630 10452 13636 10464
rect 13587 10424 13636 10452
rect 13587 10421 13599 10424
rect 13541 10415 13599 10421
rect 13630 10412 13636 10424
rect 13688 10452 13694 10464
rect 13924 10452 13952 10619
rect 13998 10616 14004 10668
rect 14056 10616 14062 10668
rect 14277 10659 14335 10665
rect 14277 10625 14289 10659
rect 14323 10656 14335 10659
rect 14642 10656 14648 10668
rect 14323 10628 14648 10656
rect 14323 10625 14335 10628
rect 14277 10619 14335 10625
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 15120 10665 15148 10696
rect 15194 10684 15200 10696
rect 15252 10724 15258 10736
rect 15930 10724 15936 10736
rect 15252 10696 15936 10724
rect 15252 10684 15258 10696
rect 15930 10684 15936 10696
rect 15988 10684 15994 10736
rect 16298 10684 16304 10736
rect 16356 10724 16362 10736
rect 16482 10724 16488 10736
rect 16356 10696 16488 10724
rect 16356 10684 16362 10696
rect 16482 10684 16488 10696
rect 16540 10684 16546 10736
rect 16592 10724 16620 10764
rect 16850 10752 16856 10804
rect 16908 10752 16914 10804
rect 17218 10724 17224 10736
rect 16592 10696 17224 10724
rect 17218 10684 17224 10696
rect 17276 10684 17282 10736
rect 17310 10684 17316 10736
rect 17368 10684 17374 10736
rect 15105 10659 15163 10665
rect 15105 10625 15117 10659
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15289 10659 15347 10665
rect 15289 10625 15301 10659
rect 15335 10656 15347 10659
rect 15378 10656 15384 10668
rect 15335 10628 15384 10656
rect 15335 10625 15347 10628
rect 15289 10619 15347 10625
rect 15378 10616 15384 10628
rect 15436 10656 15442 10668
rect 15473 10659 15531 10665
rect 15473 10656 15485 10659
rect 15436 10628 15485 10656
rect 15436 10616 15442 10628
rect 15473 10625 15485 10628
rect 15519 10625 15531 10659
rect 15473 10619 15531 10625
rect 15654 10616 15660 10668
rect 15712 10656 15718 10668
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15712 10628 15853 10656
rect 15712 10616 15718 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 16114 10616 16120 10668
rect 16172 10616 16178 10668
rect 16390 10616 16396 10668
rect 16448 10616 16454 10668
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17328 10656 17356 10684
rect 17865 10659 17923 10665
rect 17083 10628 17816 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 15565 10591 15623 10597
rect 15565 10557 15577 10591
rect 15611 10588 15623 10591
rect 15933 10591 15991 10597
rect 15933 10588 15945 10591
rect 15611 10560 15945 10588
rect 15611 10557 15623 10560
rect 15565 10551 15623 10557
rect 15933 10557 15945 10560
rect 15979 10557 15991 10591
rect 15933 10551 15991 10557
rect 17126 10548 17132 10600
rect 17184 10548 17190 10600
rect 17218 10548 17224 10600
rect 17276 10548 17282 10600
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10588 17371 10591
rect 17586 10588 17592 10600
rect 17359 10560 17592 10588
rect 17359 10557 17371 10560
rect 17313 10551 17371 10557
rect 17586 10548 17592 10560
rect 17644 10548 17650 10600
rect 17788 10597 17816 10628
rect 17865 10625 17877 10659
rect 17911 10656 17923 10659
rect 18322 10656 18328 10668
rect 17911 10628 18328 10656
rect 17911 10625 17923 10628
rect 17865 10619 17923 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 17773 10591 17831 10597
rect 17773 10557 17785 10591
rect 17819 10557 17831 10591
rect 17773 10551 17831 10557
rect 14185 10523 14243 10529
rect 14185 10489 14197 10523
rect 14231 10520 14243 10523
rect 15378 10520 15384 10532
rect 14231 10492 15384 10520
rect 14231 10489 14243 10492
rect 14185 10483 14243 10489
rect 15378 10480 15384 10492
rect 15436 10480 15442 10532
rect 15654 10480 15660 10532
rect 15712 10520 15718 10532
rect 15749 10523 15807 10529
rect 15749 10520 15761 10523
rect 15712 10492 15761 10520
rect 15712 10480 15718 10492
rect 15749 10489 15761 10492
rect 15795 10520 15807 10523
rect 17497 10523 17555 10529
rect 17497 10520 17509 10523
rect 15795 10492 17509 10520
rect 15795 10489 15807 10492
rect 15749 10483 15807 10489
rect 17497 10489 17509 10492
rect 17543 10489 17555 10523
rect 17497 10483 17555 10489
rect 13688 10424 13952 10452
rect 13688 10412 13694 10424
rect 15194 10412 15200 10464
rect 15252 10412 15258 10464
rect 15473 10455 15531 10461
rect 15473 10421 15485 10455
rect 15519 10452 15531 10455
rect 16298 10452 16304 10464
rect 15519 10424 16304 10452
rect 15519 10421 15531 10424
rect 15473 10415 15531 10421
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 17126 10412 17132 10464
rect 17184 10452 17190 10464
rect 18233 10455 18291 10461
rect 18233 10452 18245 10455
rect 17184 10424 18245 10452
rect 17184 10412 17190 10424
rect 18233 10421 18245 10424
rect 18279 10421 18291 10455
rect 18233 10415 18291 10421
rect 1104 10362 18860 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 18860 10362
rect 1104 10288 18860 10310
rect 2682 10208 2688 10260
rect 2740 10208 2746 10260
rect 5350 10248 5356 10260
rect 5184 10220 5356 10248
rect 1854 10072 1860 10124
rect 1912 10112 1918 10124
rect 2501 10115 2559 10121
rect 2501 10112 2513 10115
rect 1912 10084 2513 10112
rect 1912 10072 1918 10084
rect 2501 10081 2513 10084
rect 2547 10112 2559 10115
rect 2590 10112 2596 10124
rect 2547 10084 2596 10112
rect 2547 10081 2559 10084
rect 2501 10075 2559 10081
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1946 10044 1952 10056
rect 1596 10016 1952 10044
rect 1596 9917 1624 10016
rect 1946 10004 1952 10016
rect 2004 10044 2010 10056
rect 2774 10044 2780 10056
rect 2004 10016 2780 10044
rect 2004 10004 2010 10016
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 4706 10004 4712 10056
rect 4764 10004 4770 10056
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10044 5135 10047
rect 5184 10044 5212 10220
rect 5350 10208 5356 10220
rect 5408 10248 5414 10260
rect 5408 10220 6684 10248
rect 5408 10208 5414 10220
rect 5445 10183 5503 10189
rect 5445 10149 5457 10183
rect 5491 10149 5503 10183
rect 5445 10143 5503 10149
rect 5123 10016 5212 10044
rect 5261 10047 5319 10053
rect 5123 10013 5135 10016
rect 5077 10007 5135 10013
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5460 10044 5488 10143
rect 5307 10016 5488 10044
rect 5905 10047 5963 10053
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 4724 9976 4752 10004
rect 5920 9976 5948 10007
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6549 10047 6607 10053
rect 6549 10044 6561 10047
rect 6144 10016 6561 10044
rect 6144 10004 6150 10016
rect 6549 10013 6561 10016
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 4724 9948 6132 9976
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9877 1639 9911
rect 1581 9871 1639 9877
rect 1670 9868 1676 9920
rect 1728 9908 1734 9920
rect 2041 9911 2099 9917
rect 2041 9908 2053 9911
rect 1728 9880 2053 9908
rect 1728 9868 1734 9880
rect 2041 9877 2053 9880
rect 2087 9877 2099 9911
rect 2041 9871 2099 9877
rect 4249 9911 4307 9917
rect 4249 9877 4261 9911
rect 4295 9908 4307 9911
rect 4614 9908 4620 9920
rect 4295 9880 4620 9908
rect 4295 9877 4307 9880
rect 4249 9871 4307 9877
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9908 5319 9911
rect 5994 9908 6000 9920
rect 5307 9880 6000 9908
rect 5307 9877 5319 9880
rect 5261 9871 5319 9877
rect 5994 9868 6000 9880
rect 6052 9868 6058 9920
rect 6104 9917 6132 9948
rect 6089 9911 6147 9917
rect 6089 9877 6101 9911
rect 6135 9877 6147 9911
rect 6564 9908 6592 10007
rect 6656 9985 6684 10220
rect 7742 10208 7748 10260
rect 7800 10248 7806 10260
rect 9033 10251 9091 10257
rect 9033 10248 9045 10251
rect 7800 10220 9045 10248
rect 7800 10208 7806 10220
rect 9033 10217 9045 10220
rect 9079 10217 9091 10251
rect 9033 10211 9091 10217
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9750 10251 9808 10257
rect 9750 10248 9762 10251
rect 9548 10220 9762 10248
rect 9548 10208 9554 10220
rect 9750 10217 9762 10220
rect 9796 10217 9808 10251
rect 9750 10211 9808 10217
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10192 10220 10824 10248
rect 10192 10208 10198 10220
rect 10796 10180 10824 10220
rect 11146 10208 11152 10260
rect 11204 10248 11210 10260
rect 11241 10251 11299 10257
rect 11241 10248 11253 10251
rect 11204 10220 11253 10248
rect 11204 10208 11210 10220
rect 11241 10217 11253 10220
rect 11287 10217 11299 10251
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 11241 10211 11299 10217
rect 12406 10220 12909 10248
rect 12406 10180 12434 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 12897 10211 12955 10217
rect 13354 10208 13360 10260
rect 13412 10208 13418 10260
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 15470 10248 15476 10260
rect 15059 10220 15476 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 15470 10208 15476 10220
rect 15528 10208 15534 10260
rect 16206 10208 16212 10260
rect 16264 10208 16270 10260
rect 16298 10208 16304 10260
rect 16356 10208 16362 10260
rect 16390 10208 16396 10260
rect 16448 10248 16454 10260
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 16448 10220 16865 10248
rect 16448 10208 16454 10220
rect 16853 10217 16865 10220
rect 16899 10217 16911 10251
rect 16853 10211 16911 10217
rect 17957 10251 18015 10257
rect 17957 10217 17969 10251
rect 18003 10248 18015 10251
rect 18322 10248 18328 10260
rect 18003 10220 18328 10248
rect 18003 10217 18015 10220
rect 17957 10211 18015 10217
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 13078 10180 13084 10192
rect 10796 10152 12434 10180
rect 12820 10152 13084 10180
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10112 9551 10115
rect 9766 10112 9772 10124
rect 9539 10084 9772 10112
rect 9539 10081 9551 10084
rect 9493 10075 9551 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 12820 10121 12848 10152
rect 13078 10140 13084 10152
rect 13136 10140 13142 10192
rect 13173 10183 13231 10189
rect 13173 10149 13185 10183
rect 13219 10149 13231 10183
rect 13173 10143 13231 10149
rect 15197 10183 15255 10189
rect 15197 10149 15209 10183
rect 15243 10180 15255 10183
rect 16316 10180 16344 10208
rect 15243 10152 16344 10180
rect 15243 10149 15255 10152
rect 15197 10143 15255 10149
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10081 12863 10115
rect 12805 10075 12863 10081
rect 8021 10047 8079 10053
rect 8021 10044 8033 10047
rect 6840 10016 8033 10044
rect 6840 9985 6868 10016
rect 8021 10013 8033 10016
rect 8067 10044 8079 10047
rect 8110 10044 8116 10056
rect 8067 10016 8116 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8662 10004 8668 10056
rect 8720 10004 8726 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 6641 9979 6699 9985
rect 6641 9945 6653 9979
rect 6687 9945 6699 9979
rect 6641 9939 6699 9945
rect 6825 9979 6883 9985
rect 6825 9945 6837 9979
rect 6871 9945 6883 9979
rect 6825 9939 6883 9945
rect 6840 9908 6868 9939
rect 7374 9936 7380 9988
rect 7432 9976 7438 9988
rect 7469 9979 7527 9985
rect 7469 9976 7481 9979
rect 7432 9948 7481 9976
rect 7432 9936 7438 9948
rect 7469 9945 7481 9948
rect 7515 9945 7527 9979
rect 7469 9939 7527 9945
rect 8389 9979 8447 9985
rect 8389 9945 8401 9979
rect 8435 9976 8447 9979
rect 8570 9976 8576 9988
rect 8435 9948 8576 9976
rect 8435 9945 8447 9948
rect 8389 9939 8447 9945
rect 8570 9936 8576 9948
rect 8628 9976 8634 9988
rect 9140 9976 9168 10007
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 11517 10047 11575 10053
rect 11517 10044 11529 10047
rect 11296 10016 11529 10044
rect 11296 10004 11302 10016
rect 11517 10013 11529 10016
rect 11563 10013 11575 10047
rect 11517 10007 11575 10013
rect 12986 10004 12992 10056
rect 13044 10004 13050 10056
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10044 13139 10047
rect 13188 10044 13216 10143
rect 16482 10140 16488 10192
rect 16540 10180 16546 10192
rect 17497 10183 17555 10189
rect 17497 10180 17509 10183
rect 16540 10152 17509 10180
rect 16540 10140 16546 10152
rect 17497 10149 17509 10152
rect 17543 10149 17555 10183
rect 17497 10143 17555 10149
rect 17586 10140 17592 10192
rect 17644 10180 17650 10192
rect 18233 10183 18291 10189
rect 18233 10180 18245 10183
rect 17644 10152 18245 10180
rect 17644 10140 17650 10152
rect 18233 10149 18245 10152
rect 18279 10149 18291 10183
rect 18233 10143 18291 10149
rect 14553 10115 14611 10121
rect 14553 10081 14565 10115
rect 14599 10081 14611 10115
rect 14553 10075 14611 10081
rect 13127 10016 13216 10044
rect 13127 10013 13139 10016
rect 13081 10007 13139 10013
rect 13262 10004 13268 10056
rect 13320 10044 13326 10056
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 13320 10016 13369 10044
rect 13320 10004 13326 10016
rect 13357 10013 13369 10016
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10044 13599 10047
rect 14182 10044 14188 10056
rect 13587 10016 14188 10044
rect 13587 10013 13599 10016
rect 13541 10007 13599 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 11425 9979 11483 9985
rect 11425 9976 11437 9979
rect 8628 9948 9168 9976
rect 10994 9948 11437 9976
rect 8628 9936 8634 9948
rect 11425 9945 11437 9948
rect 11471 9945 11483 9979
rect 11425 9939 11483 9945
rect 13817 9979 13875 9985
rect 13817 9945 13829 9979
rect 13863 9976 13875 9979
rect 14093 9979 14151 9985
rect 14093 9976 14105 9979
rect 13863 9948 14105 9976
rect 13863 9945 13875 9948
rect 13817 9939 13875 9945
rect 14093 9945 14105 9948
rect 14139 9945 14151 9979
rect 14093 9939 14151 9945
rect 14384 9920 14412 10007
rect 14568 9976 14596 10075
rect 15102 10072 15108 10124
rect 15160 10072 15166 10124
rect 15286 10072 15292 10124
rect 15344 10121 15350 10124
rect 15344 10115 15384 10121
rect 15372 10112 15384 10115
rect 17773 10115 17831 10121
rect 15372 10084 16344 10112
rect 15372 10081 15384 10084
rect 15344 10075 15384 10081
rect 15344 10072 15350 10075
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15565 10047 15623 10053
rect 15565 10044 15577 10047
rect 15252 10016 15577 10044
rect 15252 10004 15258 10016
rect 15565 10013 15577 10016
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 15746 10004 15752 10056
rect 15804 10004 15810 10056
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 15378 9976 15384 9988
rect 14568 9948 15384 9976
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 15473 9979 15531 9985
rect 15473 9945 15485 9979
rect 15519 9945 15531 9979
rect 15856 9976 15884 10007
rect 15930 10004 15936 10056
rect 15988 10004 15994 10056
rect 16316 10053 16344 10084
rect 17773 10081 17785 10115
rect 17819 10112 17831 10115
rect 17954 10112 17960 10124
rect 17819 10084 17960 10112
rect 17819 10081 17831 10084
rect 17773 10075 17831 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16390 10004 16396 10056
rect 16448 10004 16454 10056
rect 17037 10047 17095 10053
rect 17037 10013 17049 10047
rect 17083 10044 17095 10047
rect 17218 10044 17224 10056
rect 17083 10016 17224 10044
rect 17083 10013 17095 10016
rect 17037 10007 17095 10013
rect 17218 10004 17224 10016
rect 17276 10004 17282 10056
rect 17310 10004 17316 10056
rect 17368 10044 17374 10056
rect 18049 10047 18107 10053
rect 18049 10044 18061 10047
rect 17368 10016 18061 10044
rect 17368 10004 17374 10016
rect 18049 10013 18061 10016
rect 18095 10013 18107 10047
rect 18049 10007 18107 10013
rect 18322 10004 18328 10056
rect 18380 10004 18386 10056
rect 15856 9948 16712 9976
rect 15473 9939 15531 9945
rect 6564 9880 6868 9908
rect 6089 9871 6147 9877
rect 7006 9868 7012 9920
rect 7064 9868 7070 9920
rect 14366 9868 14372 9920
rect 14424 9908 14430 9920
rect 15102 9908 15108 9920
rect 14424 9880 15108 9908
rect 14424 9868 14430 9880
rect 15102 9868 15108 9880
rect 15160 9868 15166 9920
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15488 9908 15516 9939
rect 15252 9880 15516 9908
rect 15252 9868 15258 9880
rect 16022 9868 16028 9920
rect 16080 9908 16086 9920
rect 16390 9908 16396 9920
rect 16080 9880 16396 9908
rect 16080 9868 16086 9880
rect 16390 9868 16396 9880
rect 16448 9868 16454 9920
rect 16684 9917 16712 9948
rect 16669 9911 16727 9917
rect 16669 9877 16681 9911
rect 16715 9877 16727 9911
rect 16669 9871 16727 9877
rect 17126 9868 17132 9920
rect 17184 9908 17190 9920
rect 17221 9911 17279 9917
rect 17221 9908 17233 9911
rect 17184 9880 17233 9908
rect 17184 9868 17190 9880
rect 17221 9877 17233 9880
rect 17267 9877 17279 9911
rect 17221 9871 17279 9877
rect 1104 9818 18860 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 18860 9818
rect 1104 9744 18860 9766
rect 1946 9704 1952 9716
rect 1504 9676 1952 9704
rect 1504 9577 1532 9676
rect 1946 9664 1952 9676
rect 2004 9664 2010 9716
rect 6181 9707 6239 9713
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 6638 9704 6644 9716
rect 6227 9676 6644 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 6638 9664 6644 9676
rect 6696 9664 6702 9716
rect 10321 9707 10379 9713
rect 10321 9673 10333 9707
rect 10367 9704 10379 9707
rect 10367 9676 10548 9704
rect 10367 9673 10379 9676
rect 10321 9667 10379 9673
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 2685 9639 2743 9645
rect 1811 9608 2544 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9537 1547 9571
rect 1489 9531 1547 9537
rect 1581 9571 1639 9577
rect 1581 9537 1593 9571
rect 1627 9568 1639 9571
rect 1670 9568 1676 9580
rect 1627 9540 1676 9568
rect 1627 9537 1639 9540
rect 1581 9531 1639 9537
rect 1670 9528 1676 9540
rect 1728 9528 1734 9580
rect 1854 9528 1860 9580
rect 1912 9528 1918 9580
rect 1946 9528 1952 9580
rect 2004 9528 2010 9580
rect 2516 9577 2544 9608
rect 2685 9605 2697 9639
rect 2731 9636 2743 9639
rect 3263 9639 3321 9645
rect 3263 9636 3275 9639
rect 2731 9608 3275 9636
rect 2731 9605 2743 9608
rect 2685 9599 2743 9605
rect 3252 9605 3275 9608
rect 3309 9605 3321 9639
rect 4706 9636 4712 9648
rect 3252 9599 3321 9605
rect 3436 9608 4712 9636
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9537 2559 9571
rect 2501 9531 2559 9537
rect 1765 9503 1823 9509
rect 1765 9469 1777 9503
rect 1811 9469 1823 9503
rect 2317 9503 2375 9509
rect 2317 9500 2329 9503
rect 1765 9463 1823 9469
rect 2240 9472 2329 9500
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 1780 9432 1808 9463
rect 2240 9444 2268 9472
rect 2317 9469 2329 9472
rect 2363 9469 2375 9503
rect 2317 9463 2375 9469
rect 2869 9503 2927 9509
rect 2869 9469 2881 9503
rect 2915 9500 2927 9503
rect 2958 9500 2964 9512
rect 2915 9472 2964 9500
rect 2915 9469 2927 9472
rect 2869 9463 2927 9469
rect 2958 9460 2964 9472
rect 3016 9460 3022 9512
rect 1636 9404 1900 9432
rect 1636 9392 1642 9404
rect 1872 9373 1900 9404
rect 2222 9392 2228 9444
rect 2280 9392 2286 9444
rect 1857 9367 1915 9373
rect 1857 9333 1869 9367
rect 1903 9364 1915 9367
rect 2314 9364 2320 9376
rect 1903 9336 2320 9364
rect 1903 9333 1915 9336
rect 1857 9327 1915 9333
rect 2314 9324 2320 9336
rect 2372 9324 2378 9376
rect 2961 9367 3019 9373
rect 2961 9333 2973 9367
rect 3007 9364 3019 9367
rect 3142 9364 3148 9376
rect 3007 9336 3148 9364
rect 3007 9333 3019 9336
rect 2961 9327 3019 9333
rect 3142 9324 3148 9336
rect 3200 9324 3206 9376
rect 3252 9364 3280 9599
rect 3436 9577 3464 9608
rect 3388 9571 3464 9577
rect 3388 9537 3400 9571
rect 3434 9540 3464 9571
rect 3605 9571 3663 9577
rect 3605 9568 3617 9571
rect 3528 9540 3617 9568
rect 3434 9537 3446 9540
rect 3388 9531 3446 9537
rect 3528 9441 3556 9540
rect 3605 9537 3617 9540
rect 3651 9537 3663 9571
rect 3605 9531 3663 9537
rect 3789 9571 3847 9577
rect 3789 9537 3801 9571
rect 3835 9568 3847 9571
rect 4062 9568 4068 9580
rect 3835 9540 4068 9568
rect 3835 9537 3847 9540
rect 3789 9531 3847 9537
rect 4062 9528 4068 9540
rect 4120 9528 4126 9580
rect 4172 9577 4200 9608
rect 4706 9596 4712 9608
rect 4764 9596 4770 9648
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 5813 9639 5871 9645
rect 5813 9636 5825 9639
rect 5684 9608 5825 9636
rect 5684 9596 5690 9608
rect 5813 9605 5825 9608
rect 5859 9605 5871 9639
rect 5813 9599 5871 9605
rect 6029 9639 6087 9645
rect 6029 9605 6041 9639
rect 6075 9636 6087 9639
rect 7006 9636 7012 9648
rect 6075 9608 7012 9636
rect 6075 9605 6087 9608
rect 6029 9599 6087 9605
rect 7006 9596 7012 9608
rect 7064 9596 7070 9648
rect 9674 9596 9680 9648
rect 9732 9636 9738 9648
rect 10410 9636 10416 9648
rect 9732 9608 10416 9636
rect 9732 9596 9738 9608
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 10520 9636 10548 9676
rect 12176 9676 13124 9704
rect 10613 9639 10671 9645
rect 10613 9636 10625 9639
rect 10520 9608 10625 9636
rect 10613 9605 10625 9608
rect 10659 9605 10671 9639
rect 10613 9599 10671 9605
rect 11057 9639 11115 9645
rect 11057 9605 11069 9639
rect 11103 9636 11115 9639
rect 12176 9636 12204 9676
rect 11103 9608 12204 9636
rect 11103 9605 11115 9608
rect 11057 9599 11115 9605
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10321 9571 10379 9577
rect 10321 9537 10333 9571
rect 10367 9568 10379 9571
rect 10962 9568 10968 9580
rect 10367 9540 10968 9568
rect 10367 9537 10379 9540
rect 10321 9531 10379 9537
rect 10962 9528 10968 9540
rect 11020 9568 11026 9580
rect 11072 9568 11100 9599
rect 12250 9596 12256 9648
rect 12308 9596 12314 9648
rect 13096 9636 13124 9676
rect 13630 9664 13636 9716
rect 13688 9664 13694 9716
rect 13906 9664 13912 9716
rect 13964 9704 13970 9716
rect 14642 9704 14648 9716
rect 13964 9676 14648 9704
rect 13964 9664 13970 9676
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 15197 9707 15255 9713
rect 15197 9673 15209 9707
rect 15243 9704 15255 9707
rect 15286 9704 15292 9716
rect 15243 9676 15292 9704
rect 15243 9673 15255 9676
rect 15197 9667 15255 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 15746 9664 15752 9716
rect 15804 9704 15810 9716
rect 15841 9707 15899 9713
rect 15841 9704 15853 9707
rect 15804 9676 15853 9704
rect 15804 9664 15810 9676
rect 15841 9673 15853 9676
rect 15887 9673 15899 9707
rect 15841 9667 15899 9673
rect 18322 9664 18328 9716
rect 18380 9664 18386 9716
rect 13541 9639 13599 9645
rect 13541 9636 13553 9639
rect 13096 9608 13553 9636
rect 13541 9605 13553 9608
rect 13587 9636 13599 9639
rect 15562 9636 15568 9648
rect 13587 9608 15568 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 11020 9540 11100 9568
rect 11020 9528 11026 9540
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 13832 9577 13860 9608
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 17218 9596 17224 9648
rect 17276 9636 17282 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 17276 9608 18245 9636
rect 17276 9596 17282 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 11241 9571 11299 9577
rect 11241 9568 11253 9571
rect 11204 9540 11253 9568
rect 11204 9528 11210 9540
rect 11241 9537 11253 9540
rect 11287 9537 11299 9571
rect 11241 9531 11299 9537
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9537 13875 9571
rect 13817 9531 13875 9537
rect 13906 9528 13912 9580
rect 13964 9528 13970 9580
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9537 14059 9571
rect 14001 9531 14059 9537
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9568 14243 9571
rect 14366 9568 14372 9580
rect 14231 9540 14372 9568
rect 14231 9537 14243 9540
rect 14185 9531 14243 9537
rect 3878 9460 3884 9512
rect 3936 9460 3942 9512
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9469 4031 9503
rect 3973 9463 4031 9469
rect 3513 9435 3571 9441
rect 3513 9401 3525 9435
rect 3559 9401 3571 9435
rect 3513 9395 3571 9401
rect 3988 9376 4016 9463
rect 9766 9460 9772 9512
rect 9824 9500 9830 9512
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 9824 9472 11529 9500
rect 9824 9460 9830 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11793 9503 11851 9509
rect 11793 9500 11805 9503
rect 11517 9463 11575 9469
rect 11624 9472 11805 9500
rect 10873 9435 10931 9441
rect 10873 9432 10885 9435
rect 10612 9404 10885 9432
rect 3970 9364 3976 9376
rect 3252 9336 3976 9364
rect 3970 9324 3976 9336
rect 4028 9324 4034 9376
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4706 9364 4712 9376
rect 4387 9336 4712 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 5994 9324 6000 9376
rect 6052 9324 6058 9376
rect 10612 9373 10640 9404
rect 10873 9401 10885 9404
rect 10919 9401 10931 9435
rect 11624 9432 11652 9472
rect 11793 9469 11805 9472
rect 11839 9469 11851 9503
rect 14016 9500 14044 9531
rect 14366 9528 14372 9540
rect 14424 9528 14430 9580
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 15289 9571 15347 9577
rect 15289 9568 15301 9571
rect 14967 9540 15301 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 15289 9537 15301 9540
rect 15335 9537 15347 9571
rect 15289 9531 15347 9537
rect 14274 9500 14280 9512
rect 11793 9463 11851 9469
rect 13832 9472 14280 9500
rect 13832 9444 13860 9472
rect 14274 9460 14280 9472
rect 14332 9500 14338 9512
rect 14936 9500 14964 9531
rect 15470 9528 15476 9580
rect 15528 9528 15534 9580
rect 15654 9568 15660 9580
rect 15712 9577 15718 9580
rect 15620 9540 15660 9568
rect 15654 9528 15660 9540
rect 15712 9531 15720 9577
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 15764 9540 16221 9568
rect 15712 9528 15718 9531
rect 14332 9472 14964 9500
rect 15197 9503 15255 9509
rect 14332 9460 14338 9472
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15381 9503 15439 9509
rect 15381 9500 15393 9503
rect 15243 9472 15393 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15381 9469 15393 9472
rect 15427 9500 15439 9503
rect 15764 9500 15792 9540
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 17954 9528 17960 9580
rect 18012 9528 18018 9580
rect 18506 9528 18512 9580
rect 18564 9528 18570 9580
rect 15427 9472 15792 9500
rect 15427 9469 15439 9472
rect 15381 9463 15439 9469
rect 16022 9460 16028 9512
rect 16080 9500 16086 9512
rect 16117 9503 16175 9509
rect 16117 9500 16129 9503
rect 16080 9472 16129 9500
rect 16080 9460 16086 9472
rect 16117 9469 16129 9472
rect 16163 9469 16175 9503
rect 16117 9463 16175 9469
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 10873 9395 10931 9401
rect 11348 9404 11652 9432
rect 10597 9367 10655 9373
rect 10597 9333 10609 9367
rect 10643 9333 10655 9367
rect 10597 9327 10655 9333
rect 10781 9367 10839 9373
rect 10781 9333 10793 9367
rect 10827 9364 10839 9367
rect 11348 9364 11376 9404
rect 13814 9392 13820 9444
rect 13872 9392 13878 9444
rect 15013 9435 15071 9441
rect 15013 9401 15025 9435
rect 15059 9432 15071 9435
rect 15470 9432 15476 9444
rect 15059 9404 15476 9432
rect 15059 9401 15071 9404
rect 15013 9395 15071 9401
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 17402 9392 17408 9444
rect 17460 9432 17466 9444
rect 17773 9435 17831 9441
rect 17773 9432 17785 9435
rect 17460 9404 17785 9432
rect 17460 9392 17466 9404
rect 17773 9401 17785 9404
rect 17819 9401 17831 9435
rect 17773 9395 17831 9401
rect 10827 9336 11376 9364
rect 16209 9367 16267 9373
rect 10827 9333 10839 9336
rect 10781 9327 10839 9333
rect 16209 9333 16221 9367
rect 16255 9364 16267 9367
rect 16298 9364 16304 9376
rect 16255 9336 16304 9364
rect 16255 9333 16267 9336
rect 16209 9327 16267 9333
rect 16298 9324 16304 9336
rect 16356 9324 16362 9376
rect 18230 9324 18236 9376
rect 18288 9324 18294 9376
rect 1104 9274 18860 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 18860 9274
rect 1104 9200 18860 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 3053 9163 3111 9169
rect 3053 9160 3065 9163
rect 1627 9132 3065 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1688 8965 1716 9132
rect 3053 9129 3065 9132
rect 3099 9160 3111 9163
rect 3326 9160 3332 9172
rect 3099 9132 3332 9160
rect 3099 9129 3111 9132
rect 3053 9123 3111 9129
rect 3326 9120 3332 9132
rect 3384 9120 3390 9172
rect 3878 9120 3884 9172
rect 3936 9160 3942 9172
rect 4893 9163 4951 9169
rect 3936 9132 4844 9160
rect 3936 9120 3942 9132
rect 2501 9095 2559 9101
rect 2501 9061 2513 9095
rect 2547 9092 2559 9095
rect 2958 9092 2964 9104
rect 2547 9064 2964 9092
rect 2547 9061 2559 9064
rect 2501 9055 2559 9061
rect 2958 9052 2964 9064
rect 3016 9092 3022 9104
rect 4709 9095 4767 9101
rect 3016 9064 3280 9092
rect 3016 9052 3022 9064
rect 2222 8984 2228 9036
rect 2280 8984 2286 9036
rect 2314 8984 2320 9036
rect 2372 9024 2378 9036
rect 2869 9027 2927 9033
rect 2869 9024 2881 9027
rect 2372 8996 2881 9024
rect 2372 8984 2378 8996
rect 2869 8993 2881 8996
rect 2915 8993 2927 9027
rect 2869 8987 2927 8993
rect 3252 9024 3280 9064
rect 4709 9061 4721 9095
rect 4755 9061 4767 9095
rect 4816 9092 4844 9132
rect 4893 9129 4905 9163
rect 4939 9160 4951 9163
rect 5442 9160 5448 9172
rect 4939 9132 5448 9160
rect 4939 9129 4951 9132
rect 4893 9123 4951 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8904 9132 8953 9160
rect 8904 9120 8910 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 10134 9120 10140 9172
rect 10192 9160 10198 9172
rect 10686 9160 10692 9172
rect 10192 9132 10692 9160
rect 10192 9120 10198 9132
rect 10686 9120 10692 9132
rect 10744 9160 10750 9172
rect 10962 9160 10968 9172
rect 10744 9132 10968 9160
rect 10744 9120 10750 9132
rect 10962 9120 10968 9132
rect 11020 9120 11026 9172
rect 11977 9163 12035 9169
rect 11977 9129 11989 9163
rect 12023 9160 12035 9163
rect 12250 9160 12256 9172
rect 12023 9132 12256 9160
rect 12023 9129 12035 9132
rect 11977 9123 12035 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 15470 9120 15476 9172
rect 15528 9160 15534 9172
rect 16761 9163 16819 9169
rect 16761 9160 16773 9163
rect 15528 9132 16773 9160
rect 15528 9120 15534 9132
rect 16761 9129 16773 9132
rect 16807 9129 16819 9163
rect 17310 9160 17316 9172
rect 16761 9123 16819 9129
rect 16960 9132 17316 9160
rect 5074 9092 5080 9104
rect 4816 9064 5080 9092
rect 4709 9055 4767 9061
rect 3510 9024 3516 9036
rect 3252 8996 3516 9024
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2130 8956 2136 8968
rect 1811 8928 2136 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 2130 8916 2136 8928
rect 2188 8916 2194 8968
rect 2774 8916 2780 8968
rect 2832 8916 2838 8968
rect 3252 8965 3280 8996
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 3605 9027 3663 9033
rect 3605 8993 3617 9027
rect 3651 9024 3663 9027
rect 4065 9027 4123 9033
rect 4065 9024 4077 9027
rect 3651 8996 4077 9024
rect 3651 8993 3663 8996
rect 3605 8987 3663 8993
rect 4065 8993 4077 8996
rect 4111 8993 4123 9027
rect 4065 8987 4123 8993
rect 4157 9027 4215 9033
rect 4157 8993 4169 9027
rect 4203 9024 4215 9027
rect 4614 9024 4620 9036
rect 4203 8996 4620 9024
rect 4203 8993 4215 8996
rect 4157 8987 4215 8993
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4724 9024 4752 9055
rect 5074 9052 5080 9064
rect 5132 9092 5138 9104
rect 5721 9095 5779 9101
rect 5721 9092 5733 9095
rect 5132 9064 5733 9092
rect 5132 9052 5138 9064
rect 5721 9061 5733 9064
rect 5767 9061 5779 9095
rect 5721 9055 5779 9061
rect 8297 9095 8355 9101
rect 8297 9061 8309 9095
rect 8343 9092 8355 9095
rect 8665 9095 8723 9101
rect 8343 9064 8616 9092
rect 8343 9061 8355 9064
rect 8297 9055 8355 9061
rect 4890 9024 4896 9036
rect 4724 8996 4896 9024
rect 4890 8984 4896 8996
rect 4948 8984 4954 9036
rect 5813 9027 5871 9033
rect 5813 9024 5825 9027
rect 5000 8996 5825 9024
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 3786 8956 3792 8968
rect 3467 8928 3792 8956
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 3050 8848 3056 8900
rect 3108 8848 3114 8900
rect 3142 8848 3148 8900
rect 3200 8888 3206 8900
rect 3436 8888 3464 8919
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 3970 8916 3976 8968
rect 4028 8916 4034 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4338 8956 4344 8968
rect 4295 8928 4344 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4338 8916 4344 8928
rect 4396 8956 4402 8968
rect 4798 8956 4804 8968
rect 4396 8928 4804 8956
rect 4396 8916 4402 8928
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 3200 8860 3464 8888
rect 3200 8848 3206 8860
rect 2590 8780 2596 8832
rect 2648 8780 2654 8832
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 3970 8820 3976 8832
rect 3835 8792 3976 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4877 8823 4935 8829
rect 4877 8789 4889 8823
rect 4923 8820 4935 8823
rect 5000 8820 5028 8996
rect 5368 8965 5396 8996
rect 5813 8993 5825 8996
rect 5859 8993 5871 9027
rect 8018 9024 8024 9036
rect 5813 8987 5871 8993
rect 7116 8996 8024 9024
rect 5169 8959 5227 8965
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5353 8959 5411 8965
rect 5215 8928 5304 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5074 8848 5080 8900
rect 5132 8848 5138 8900
rect 4923 8792 5028 8820
rect 5276 8820 5304 8928
rect 5353 8925 5365 8959
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8956 6055 8959
rect 6086 8956 6092 8968
rect 6043 8928 6092 8956
rect 6043 8925 6055 8928
rect 5997 8919 6055 8925
rect 6086 8916 6092 8928
rect 6144 8916 6150 8968
rect 6178 8916 6184 8968
rect 6236 8916 6242 8968
rect 7116 8965 7144 8996
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 8386 8984 8392 9036
rect 8444 8984 8450 9036
rect 8588 9024 8616 9064
rect 8665 9061 8677 9095
rect 8711 9092 8723 9095
rect 9122 9092 9128 9104
rect 8711 9064 9128 9092
rect 8711 9061 8723 9064
rect 8665 9055 8723 9061
rect 9122 9052 9128 9064
rect 9180 9052 9186 9104
rect 9030 9024 9036 9036
rect 8588 8996 9036 9024
rect 9030 8984 9036 8996
rect 9088 9024 9094 9036
rect 9490 9024 9496 9036
rect 9088 8996 9496 9024
rect 9088 8984 9094 8996
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10652 8996 10701 9024
rect 10652 8984 10658 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 7101 8959 7159 8965
rect 7101 8925 7113 8959
rect 7147 8925 7159 8959
rect 7101 8919 7159 8925
rect 7194 8959 7252 8965
rect 7194 8925 7206 8959
rect 7240 8925 7252 8959
rect 7194 8919 7252 8925
rect 5442 8848 5448 8900
rect 5500 8848 5506 8900
rect 6270 8848 6276 8900
rect 6328 8888 6334 8900
rect 7209 8888 7237 8919
rect 7374 8916 7380 8968
rect 7432 8916 7438 8968
rect 7566 8959 7624 8965
rect 7566 8925 7578 8959
rect 7612 8925 7624 8959
rect 7566 8919 7624 8925
rect 8168 8959 8226 8965
rect 8168 8925 8180 8959
rect 8214 8956 8226 8959
rect 8294 8956 8300 8968
rect 8214 8928 8300 8956
rect 8214 8925 8226 8928
rect 8168 8919 8226 8925
rect 6328 8860 7237 8888
rect 6328 8848 6334 8860
rect 7282 8848 7288 8900
rect 7340 8888 7346 8900
rect 7469 8891 7527 8897
rect 7469 8888 7481 8891
rect 7340 8860 7481 8888
rect 7340 8848 7346 8860
rect 7469 8857 7481 8860
rect 7515 8857 7527 8891
rect 7469 8851 7527 8857
rect 5350 8820 5356 8832
rect 5276 8792 5356 8820
rect 4923 8789 4935 8792
rect 4877 8783 4935 8789
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5534 8780 5540 8832
rect 5592 8780 5598 8832
rect 7190 8780 7196 8832
rect 7248 8820 7254 8832
rect 7576 8820 7604 8919
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 8021 8891 8079 8897
rect 8021 8857 8033 8891
rect 8067 8857 8079 8891
rect 9140 8888 9168 8919
rect 9306 8916 9312 8968
rect 9364 8916 9370 8968
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 10413 8959 10471 8965
rect 10413 8925 10425 8959
rect 10459 8956 10471 8959
rect 10459 8928 11192 8956
rect 10459 8925 10471 8928
rect 10413 8919 10471 8925
rect 9214 8888 9220 8900
rect 9140 8860 9220 8888
rect 8021 8851 8079 8857
rect 7248 8792 7604 8820
rect 7745 8823 7803 8829
rect 7248 8780 7254 8792
rect 7745 8789 7757 8823
rect 7791 8820 7803 8823
rect 8036 8820 8064 8851
rect 9214 8848 9220 8860
rect 9272 8888 9278 8900
rect 10134 8888 10140 8900
rect 9272 8860 10140 8888
rect 9272 8848 9278 8860
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 11164 8888 11192 8928
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11296 8928 11897 8956
rect 11296 8916 11302 8928
rect 11885 8925 11897 8928
rect 11931 8956 11943 8959
rect 12158 8956 12164 8968
rect 11931 8928 12164 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 16850 8956 16856 8968
rect 16807 8928 16856 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 16960 8965 16988 9132
rect 17310 9120 17316 9132
rect 17368 9160 17374 9172
rect 17865 9163 17923 9169
rect 17865 9160 17877 9163
rect 17368 9132 17877 9160
rect 17368 9120 17374 9132
rect 17865 9129 17877 9132
rect 17911 9129 17923 9163
rect 17865 9123 17923 9129
rect 17957 9163 18015 9169
rect 17957 9129 17969 9163
rect 18003 9160 18015 9163
rect 18046 9160 18052 9172
rect 18003 9132 18052 9160
rect 18003 9129 18015 9132
rect 17957 9123 18015 9129
rect 18046 9120 18052 9132
rect 18104 9120 18110 9172
rect 18417 9163 18475 9169
rect 18417 9129 18429 9163
rect 18463 9160 18475 9163
rect 18506 9160 18512 9172
rect 18463 9132 18512 9160
rect 18463 9129 18475 9132
rect 18417 9123 18475 9129
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 17218 8984 17224 9036
rect 17276 8984 17282 9036
rect 18322 9024 18328 9036
rect 18156 8996 18328 9024
rect 16945 8959 17003 8965
rect 16945 8925 16957 8959
rect 16991 8925 17003 8959
rect 16945 8919 17003 8925
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 18156 8965 18184 8996
rect 18322 8984 18328 8996
rect 18380 8984 18386 9036
rect 18141 8959 18199 8965
rect 17460 8928 18092 8956
rect 17460 8916 17466 8928
rect 18064 8900 18092 8928
rect 18141 8925 18153 8959
rect 18187 8925 18199 8959
rect 18141 8919 18199 8925
rect 18230 8916 18236 8968
rect 18288 8916 18294 8968
rect 11330 8888 11336 8900
rect 11164 8860 11336 8888
rect 11330 8848 11336 8860
rect 11388 8888 11394 8900
rect 13538 8888 13544 8900
rect 11388 8860 13544 8888
rect 11388 8848 11394 8860
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 17678 8848 17684 8900
rect 17736 8897 17742 8900
rect 17736 8891 17764 8897
rect 17752 8857 17764 8891
rect 17736 8851 17764 8857
rect 17736 8848 17742 8851
rect 18046 8848 18052 8900
rect 18104 8888 18110 8900
rect 18417 8891 18475 8897
rect 18417 8888 18429 8891
rect 18104 8860 18429 8888
rect 18104 8848 18110 8860
rect 18417 8857 18429 8860
rect 18463 8857 18475 8891
rect 18417 8851 18475 8857
rect 7791 8792 8064 8820
rect 7791 8789 7803 8792
rect 7745 8783 7803 8789
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 10778 8820 10784 8832
rect 9916 8792 10784 8820
rect 9916 8780 9922 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 17218 8820 17224 8832
rect 16264 8792 17224 8820
rect 16264 8780 16270 8792
rect 17218 8780 17224 8792
rect 17276 8820 17282 8832
rect 17497 8823 17555 8829
rect 17497 8820 17509 8823
rect 17276 8792 17509 8820
rect 17276 8780 17282 8792
rect 17497 8789 17509 8792
rect 17543 8789 17555 8823
rect 17497 8783 17555 8789
rect 17586 8780 17592 8832
rect 17644 8780 17650 8832
rect 1104 8730 18860 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 18860 8730
rect 1104 8656 18860 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2372 8588 3556 8616
rect 2372 8576 2378 8588
rect 3050 8548 3056 8560
rect 2332 8520 3056 8548
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2332 8489 2360 8520
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 2317 8483 2375 8489
rect 2317 8480 2329 8483
rect 1912 8452 2329 8480
rect 1912 8440 1918 8452
rect 2317 8449 2329 8452
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 3528 8489 3556 8588
rect 4338 8576 4344 8628
rect 4396 8576 4402 8628
rect 4890 8616 4896 8628
rect 4540 8588 4896 8616
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3660 8520 3985 8548
rect 3660 8508 3666 8520
rect 3973 8517 3985 8520
rect 4019 8517 4031 8551
rect 3973 8511 4031 8517
rect 4065 8551 4123 8557
rect 4065 8517 4077 8551
rect 4111 8548 4123 8551
rect 4540 8548 4568 8588
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8616 5043 8619
rect 5166 8616 5172 8628
rect 5031 8588 5172 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 8294 8576 8300 8628
rect 8352 8576 8358 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 8772 8588 9321 8616
rect 6086 8548 6092 8560
rect 4111 8520 4568 8548
rect 4632 8520 6092 8548
rect 4111 8517 4123 8520
rect 4065 8511 4123 8517
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 4154 8440 4160 8492
rect 4212 8440 4218 8492
rect 4632 8480 4660 8520
rect 6086 8508 6092 8520
rect 6144 8548 6150 8560
rect 7469 8551 7527 8557
rect 6144 8520 7052 8548
rect 6144 8508 6150 8520
rect 4264 8452 4660 8480
rect 1394 8372 1400 8424
rect 1452 8372 1458 8424
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8412 1731 8415
rect 2516 8412 2544 8440
rect 1719 8384 2544 8412
rect 2685 8415 2743 8421
rect 1719 8381 1731 8384
rect 1673 8375 1731 8381
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 2774 8412 2780 8424
rect 2731 8384 2780 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 2774 8372 2780 8384
rect 2832 8372 2838 8424
rect 3421 8415 3479 8421
rect 3421 8381 3433 8415
rect 3467 8381 3479 8415
rect 3421 8375 3479 8381
rect 2482 8347 2540 8353
rect 2482 8313 2494 8347
rect 2528 8344 2540 8347
rect 3145 8347 3203 8353
rect 3145 8344 3157 8347
rect 2528 8316 3157 8344
rect 2528 8313 2540 8316
rect 2482 8307 2540 8313
rect 3145 8313 3157 8316
rect 3191 8313 3203 8347
rect 3145 8307 3203 8313
rect 3234 8304 3240 8356
rect 3292 8344 3298 8356
rect 3436 8344 3464 8375
rect 4264 8344 4292 8452
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8480 4859 8483
rect 5258 8480 5264 8492
rect 4847 8452 5264 8480
rect 4847 8449 4859 8452
rect 4801 8443 4859 8449
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 4522 8372 4528 8424
rect 4580 8372 4586 8424
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8381 4675 8415
rect 4617 8375 4675 8381
rect 3292 8316 4292 8344
rect 4632 8344 4660 8375
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 5736 8412 5764 8443
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8480 6055 8483
rect 6178 8480 6184 8492
rect 6043 8452 6184 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6454 8440 6460 8492
rect 6512 8440 6518 8492
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 7024 8489 7052 8520
rect 7469 8517 7481 8551
rect 7515 8548 7527 8551
rect 8018 8548 8024 8560
rect 7515 8520 8024 8548
rect 7515 8517 7527 8520
rect 7469 8511 7527 8517
rect 8018 8508 8024 8520
rect 8076 8548 8082 8560
rect 8076 8520 8708 8548
rect 8076 8508 8082 8520
rect 6917 8483 6975 8489
rect 6917 8449 6929 8483
rect 6963 8449 6975 8483
rect 6917 8443 6975 8449
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 6089 8415 6147 8421
rect 6089 8412 6101 8415
rect 5684 8384 6101 8412
rect 5684 8372 5690 8384
rect 6089 8381 6101 8384
rect 6135 8412 6147 8415
rect 6932 8412 6960 8443
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 7834 8480 7840 8492
rect 7340 8452 7840 8480
rect 7340 8440 7346 8452
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 7926 8440 7932 8492
rect 7984 8440 7990 8492
rect 8113 8483 8171 8489
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8478 8480 8484 8492
rect 8159 8452 8484 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8478 8440 8484 8452
rect 8536 8440 8542 8492
rect 6135 8384 6960 8412
rect 7101 8415 7159 8421
rect 6135 8381 6147 8384
rect 6089 8375 6147 8381
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7190 8412 7196 8424
rect 7147 8384 7196 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 4706 8344 4712 8356
rect 4632 8316 4712 8344
rect 3292 8304 3298 8316
rect 4706 8304 4712 8316
rect 4764 8304 4770 8356
rect 4890 8304 4896 8356
rect 4948 8344 4954 8356
rect 5442 8344 5448 8356
rect 4948 8316 5448 8344
rect 4948 8304 4954 8316
rect 5442 8304 5448 8316
rect 5500 8344 5506 8356
rect 6454 8344 6460 8356
rect 5500 8316 6460 8344
rect 5500 8304 5506 8316
rect 6454 8304 6460 8316
rect 6512 8304 6518 8356
rect 6549 8347 6607 8353
rect 6549 8313 6561 8347
rect 6595 8344 6607 8347
rect 7116 8344 7144 8375
rect 7190 8372 7196 8384
rect 7248 8372 7254 8424
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8260 8384 8585 8412
rect 8260 8372 8266 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8680 8412 8708 8520
rect 8772 8489 8800 8588
rect 9309 8585 9321 8588
rect 9355 8616 9367 8619
rect 9398 8616 9404 8628
rect 9355 8588 9404 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9490 8576 9496 8628
rect 9548 8616 9554 8628
rect 10597 8619 10655 8625
rect 10597 8616 10609 8619
rect 9548 8588 10609 8616
rect 9548 8576 9554 8588
rect 10597 8585 10609 8588
rect 10643 8585 10655 8619
rect 10597 8579 10655 8585
rect 12986 8576 12992 8628
rect 13044 8616 13050 8628
rect 13265 8619 13323 8625
rect 13265 8616 13277 8619
rect 13044 8588 13277 8616
rect 13044 8576 13050 8588
rect 13265 8585 13277 8588
rect 13311 8585 13323 8619
rect 13265 8579 13323 8585
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14461 8619 14519 8625
rect 14461 8616 14473 8619
rect 14056 8588 14473 8616
rect 14056 8576 14062 8588
rect 14461 8585 14473 8588
rect 14507 8585 14519 8619
rect 14461 8579 14519 8585
rect 16850 8576 16856 8628
rect 16908 8576 16914 8628
rect 17678 8576 17684 8628
rect 17736 8616 17742 8628
rect 17773 8619 17831 8625
rect 17773 8616 17785 8619
rect 17736 8588 17785 8616
rect 17736 8576 17742 8588
rect 17773 8585 17785 8588
rect 17819 8585 17831 8619
rect 18506 8616 18512 8628
rect 17773 8579 17831 8585
rect 17874 8588 18512 8616
rect 8941 8551 8999 8557
rect 8941 8517 8953 8551
rect 8987 8548 8999 8551
rect 9125 8551 9183 8557
rect 9125 8548 9137 8551
rect 8987 8520 9137 8548
rect 8987 8517 8999 8520
rect 8941 8511 8999 8517
rect 9125 8517 9137 8520
rect 9171 8517 9183 8551
rect 9125 8511 9183 8517
rect 9766 8508 9772 8560
rect 9824 8548 9830 8560
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 9824 8520 10057 8548
rect 9824 8508 9830 8520
rect 10045 8517 10057 8520
rect 10091 8517 10103 8551
rect 10045 8511 10103 8517
rect 11514 8508 11520 8560
rect 11572 8548 11578 8560
rect 11977 8551 12035 8557
rect 11977 8548 11989 8551
rect 11572 8520 11989 8548
rect 11572 8508 11578 8520
rect 11977 8517 11989 8520
rect 12023 8517 12035 8551
rect 14090 8548 14096 8560
rect 11977 8511 12035 8517
rect 13556 8520 14096 8548
rect 8772 8483 8852 8489
rect 8772 8452 8806 8483
rect 8794 8449 8806 8452
rect 8840 8449 8852 8483
rect 8794 8443 8852 8449
rect 9033 8483 9091 8489
rect 9033 8449 9045 8483
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 9048 8412 9076 8443
rect 9214 8440 9220 8492
rect 9272 8440 9278 8492
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9456 8452 9505 8480
rect 9456 8440 9462 8452
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 9493 8443 9551 8449
rect 9585 8483 9643 8489
rect 9585 8449 9597 8483
rect 9631 8449 9643 8483
rect 9585 8443 9643 8449
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9677 8443 9735 8449
rect 8680 8384 9076 8412
rect 8573 8375 8631 8381
rect 6595 8316 7144 8344
rect 8021 8347 8079 8353
rect 6595 8313 6607 8316
rect 6549 8307 6607 8313
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8938 8344 8944 8356
rect 8067 8316 8944 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8938 8304 8944 8316
rect 8996 8304 9002 8356
rect 9600 8344 9628 8443
rect 9692 8412 9720 8443
rect 9858 8440 9864 8492
rect 9916 8440 9922 8492
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 13556 8489 13584 8520
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 17874 8548 17902 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 17144 8520 17902 8548
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 13540 8483 13598 8489
rect 13540 8449 13552 8483
rect 13586 8449 13598 8483
rect 13540 8443 13598 8449
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 9950 8412 9956 8424
rect 9692 8384 9956 8412
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 10318 8412 10324 8424
rect 10100 8384 10324 8412
rect 10100 8372 10106 8384
rect 10318 8372 10324 8384
rect 10376 8412 10382 8424
rect 10704 8412 10732 8443
rect 10376 8384 10732 8412
rect 10376 8372 10382 8384
rect 11808 8344 11836 8443
rect 13262 8372 13268 8424
rect 13320 8412 13326 8424
rect 13648 8412 13676 8443
rect 13722 8440 13728 8492
rect 13780 8440 13786 8492
rect 13906 8440 13912 8492
rect 13964 8440 13970 8492
rect 14277 8483 14335 8489
rect 14277 8449 14289 8483
rect 14323 8480 14335 8483
rect 14366 8480 14372 8492
rect 14323 8452 14372 8480
rect 14323 8449 14335 8452
rect 14277 8443 14335 8449
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 17034 8480 17040 8492
rect 15528 8452 17040 8480
rect 15528 8440 15534 8452
rect 17034 8440 17040 8452
rect 17092 8480 17098 8492
rect 17144 8489 17172 8520
rect 17129 8483 17187 8489
rect 17129 8480 17141 8483
rect 17092 8452 17141 8480
rect 17092 8440 17098 8452
rect 17129 8449 17141 8452
rect 17175 8449 17187 8483
rect 17129 8443 17187 8449
rect 17313 8483 17371 8489
rect 17313 8449 17325 8483
rect 17359 8480 17371 8483
rect 17494 8480 17500 8492
rect 17359 8452 17500 8480
rect 17359 8449 17371 8452
rect 17313 8443 17371 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17874 8489 17902 8520
rect 18414 8508 18420 8560
rect 18472 8508 18478 8560
rect 17589 8483 17647 8489
rect 17589 8449 17601 8483
rect 17635 8480 17647 8483
rect 17681 8483 17739 8489
rect 17681 8480 17693 8483
rect 17635 8452 17693 8480
rect 17635 8449 17647 8452
rect 17589 8443 17647 8449
rect 17681 8449 17693 8452
rect 17727 8449 17739 8483
rect 17681 8443 17739 8449
rect 17859 8483 17917 8489
rect 17859 8449 17871 8483
rect 17905 8449 17917 8483
rect 17859 8443 17917 8449
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8480 18015 8483
rect 18046 8480 18052 8492
rect 18003 8452 18052 8480
rect 18003 8449 18015 8452
rect 17957 8443 18015 8449
rect 13320 8384 13676 8412
rect 13320 8372 13326 8384
rect 13998 8372 14004 8424
rect 14056 8372 14062 8424
rect 14093 8415 14151 8421
rect 14093 8381 14105 8415
rect 14139 8381 14151 8415
rect 17696 8412 17724 8443
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18230 8412 18236 8424
rect 17696 8384 18236 8412
rect 14093 8375 14151 8381
rect 12342 8344 12348 8356
rect 9600 8316 9720 8344
rect 11808 8316 12348 8344
rect 9692 8288 9720 8316
rect 12342 8304 12348 8316
rect 12400 8344 12406 8356
rect 13814 8344 13820 8356
rect 12400 8316 13820 8344
rect 12400 8304 12406 8316
rect 13814 8304 13820 8316
rect 13872 8344 13878 8356
rect 14108 8344 14136 8375
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 13872 8316 14136 8344
rect 17221 8347 17279 8353
rect 13872 8304 13878 8316
rect 17221 8313 17233 8347
rect 17267 8344 17279 8347
rect 17310 8344 17316 8356
rect 17267 8316 17316 8344
rect 17267 8313 17279 8316
rect 17221 8307 17279 8313
rect 17310 8304 17316 8316
rect 17368 8344 17374 8356
rect 17954 8344 17960 8356
rect 17368 8316 17960 8344
rect 17368 8304 17374 8316
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 2593 8279 2651 8285
rect 2593 8245 2605 8279
rect 2639 8276 2651 8279
rect 2682 8276 2688 8288
rect 2639 8248 2688 8276
rect 2639 8245 2651 8248
rect 2593 8239 2651 8245
rect 2682 8236 2688 8248
rect 2740 8236 2746 8288
rect 2958 8236 2964 8288
rect 3016 8236 3022 8288
rect 3326 8236 3332 8288
rect 3384 8236 3390 8288
rect 5810 8236 5816 8288
rect 5868 8236 5874 8288
rect 8665 8279 8723 8285
rect 8665 8245 8677 8279
rect 8711 8276 8723 8279
rect 9214 8276 9220 8288
rect 8711 8248 9220 8276
rect 8711 8245 8723 8248
rect 8665 8239 8723 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 9674 8236 9680 8288
rect 9732 8236 9738 8288
rect 11606 8236 11612 8288
rect 11664 8236 11670 8288
rect 17402 8236 17408 8288
rect 17460 8236 17466 8288
rect 17862 8236 17868 8288
rect 17920 8276 17926 8288
rect 18049 8279 18107 8285
rect 18049 8276 18061 8279
rect 17920 8248 18061 8276
rect 17920 8236 17926 8248
rect 18049 8245 18061 8248
rect 18095 8245 18107 8279
rect 18049 8239 18107 8245
rect 18230 8236 18236 8288
rect 18288 8276 18294 8288
rect 18325 8279 18383 8285
rect 18325 8276 18337 8279
rect 18288 8248 18337 8276
rect 18288 8236 18294 8248
rect 18325 8245 18337 8248
rect 18371 8276 18383 8279
rect 18414 8276 18420 8288
rect 18371 8248 18420 8276
rect 18371 8245 18383 8248
rect 18325 8239 18383 8245
rect 18414 8236 18420 8248
rect 18472 8236 18478 8288
rect 1104 8186 18860 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 18860 8186
rect 1104 8112 18860 8134
rect 2869 8075 2927 8081
rect 2869 8041 2881 8075
rect 2915 8072 2927 8075
rect 4062 8072 4068 8084
rect 2915 8044 4068 8072
rect 2915 8041 2927 8044
rect 2869 8035 2927 8041
rect 4062 8032 4068 8044
rect 4120 8032 4126 8084
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4614 8072 4620 8084
rect 4571 8044 4620 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 7561 8075 7619 8081
rect 7561 8041 7573 8075
rect 7607 8072 7619 8075
rect 7926 8072 7932 8084
rect 7607 8044 7932 8072
rect 7607 8041 7619 8044
rect 7561 8035 7619 8041
rect 7926 8032 7932 8044
rect 7984 8032 7990 8084
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 9217 8075 9275 8081
rect 9217 8041 9229 8075
rect 9263 8072 9275 8075
rect 9306 8072 9312 8084
rect 9263 8044 9312 8072
rect 9263 8041 9275 8044
rect 9217 8035 9275 8041
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 10134 8032 10140 8084
rect 10192 8032 10198 8084
rect 10965 8075 11023 8081
rect 10965 8041 10977 8075
rect 11011 8072 11023 8075
rect 11606 8072 11612 8084
rect 11011 8044 11612 8072
rect 11011 8041 11023 8044
rect 10965 8035 11023 8041
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 14182 8032 14188 8084
rect 14240 8032 14246 8084
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 15565 8075 15623 8081
rect 15565 8072 15577 8075
rect 14599 8044 15577 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 15565 8041 15577 8044
rect 15611 8041 15623 8075
rect 18325 8075 18383 8081
rect 18325 8072 18337 8075
rect 15565 8035 15623 8041
rect 15856 8044 18337 8072
rect 4080 8004 4108 8032
rect 6822 8004 6828 8016
rect 4080 7976 4844 8004
rect 2590 7896 2596 7948
rect 2648 7896 2654 7948
rect 2958 7896 2964 7948
rect 3016 7936 3022 7948
rect 3145 7939 3203 7945
rect 3145 7936 3157 7939
rect 3016 7908 3157 7936
rect 3016 7896 3022 7908
rect 3145 7905 3157 7908
rect 3191 7905 3203 7939
rect 4617 7939 4675 7945
rect 4617 7936 4629 7939
rect 3145 7899 3203 7905
rect 4172 7908 4629 7936
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 1688 7800 1716 7831
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 3234 7868 3240 7880
rect 2556 7840 3240 7868
rect 2556 7828 2562 7840
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 3970 7828 3976 7880
rect 4028 7828 4034 7880
rect 4172 7877 4200 7908
rect 4617 7905 4629 7908
rect 4663 7936 4675 7939
rect 4706 7936 4712 7948
rect 4663 7908 4712 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 4816 7877 4844 7976
rect 5552 7976 6828 8004
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7905 5135 7939
rect 5077 7899 5135 7905
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 2682 7800 2688 7812
rect 1688 7772 2688 7800
rect 2682 7760 2688 7772
rect 2740 7760 2746 7812
rect 4246 7760 4252 7812
rect 4304 7760 4310 7812
rect 4356 7800 4384 7831
rect 4890 7828 4896 7880
rect 4948 7828 4954 7880
rect 5092 7800 5120 7899
rect 5552 7880 5580 7976
rect 6822 7964 6828 7976
rect 6880 8004 6886 8016
rect 7285 8007 7343 8013
rect 7285 8004 7297 8007
rect 6880 7976 7297 8004
rect 6880 7964 6886 7976
rect 7285 7973 7297 7976
rect 7331 7973 7343 8007
rect 7285 7967 7343 7973
rect 8202 7964 8208 8016
rect 8260 7964 8266 8016
rect 13906 7964 13912 8016
rect 13964 8004 13970 8016
rect 14645 8007 14703 8013
rect 14645 8004 14657 8007
rect 13964 7976 14657 8004
rect 13964 7964 13970 7976
rect 14645 7973 14657 7976
rect 14691 8004 14703 8007
rect 15013 8007 15071 8013
rect 15013 8004 15025 8007
rect 14691 7976 15025 8004
rect 14691 7973 14703 7976
rect 14645 7967 14703 7973
rect 15013 7973 15025 7976
rect 15059 7973 15071 8007
rect 15013 7967 15071 7973
rect 15102 7964 15108 8016
rect 15160 7964 15166 8016
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 8220 7936 8248 7964
rect 6779 7908 8248 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7868 5227 7871
rect 5534 7868 5540 7880
rect 5215 7840 5540 7868
rect 5215 7837 5227 7840
rect 5169 7831 5227 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 6086 7868 6092 7880
rect 5767 7840 6092 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6181 7871 6239 7877
rect 6181 7837 6193 7871
rect 6227 7868 6239 7871
rect 6270 7868 6276 7880
rect 6227 7840 6276 7868
rect 6227 7837 6239 7840
rect 6181 7831 6239 7837
rect 6270 7828 6276 7840
rect 6328 7828 6334 7880
rect 6365 7871 6423 7877
rect 6365 7837 6377 7871
rect 6411 7868 6423 7871
rect 6411 7840 7144 7868
rect 6411 7837 6423 7840
rect 6365 7831 6423 7837
rect 4356 7772 5120 7800
rect 3513 7735 3571 7741
rect 3513 7701 3525 7735
rect 3559 7732 3571 7735
rect 4356 7732 4384 7772
rect 6914 7760 6920 7812
rect 6972 7800 6978 7812
rect 7009 7803 7067 7809
rect 7009 7800 7021 7803
rect 6972 7772 7021 7800
rect 6972 7760 6978 7772
rect 7009 7769 7021 7772
rect 7055 7769 7067 7803
rect 7116 7800 7144 7840
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 7944 7877 7972 7908
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10870 7936 10876 7948
rect 9824 7908 10876 7936
rect 9824 7896 9830 7908
rect 10870 7896 10876 7908
rect 10928 7936 10934 7948
rect 11241 7939 11299 7945
rect 11241 7936 11253 7939
rect 10928 7908 11253 7936
rect 10928 7896 10934 7908
rect 11241 7905 11253 7908
rect 11287 7905 11299 7939
rect 11241 7899 11299 7905
rect 12066 7896 12072 7948
rect 12124 7936 12130 7948
rect 13449 7939 13507 7945
rect 13449 7936 13461 7939
rect 12124 7908 13461 7936
rect 12124 7896 12130 7908
rect 13449 7905 13461 7908
rect 13495 7905 13507 7939
rect 13449 7899 13507 7905
rect 13541 7939 13599 7945
rect 13541 7905 13553 7939
rect 13587 7936 13599 7939
rect 14366 7936 14372 7948
rect 13587 7908 14372 7936
rect 13587 7905 13599 7908
rect 13541 7899 13599 7905
rect 7699 7871 7757 7877
rect 7699 7868 7711 7871
rect 7248 7840 7711 7868
rect 7248 7828 7254 7840
rect 7699 7837 7711 7840
rect 7745 7837 7757 7871
rect 7699 7831 7757 7837
rect 7929 7871 7987 7877
rect 7929 7837 7941 7871
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8018 7828 8024 7880
rect 8076 7877 8082 7880
rect 8076 7871 8115 7877
rect 8103 7837 8115 7871
rect 8076 7831 8115 7837
rect 8076 7828 8082 7831
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 8260 7840 8309 7868
rect 8260 7828 8266 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 8444 7840 8489 7868
rect 8444 7828 8450 7840
rect 8938 7828 8944 7880
rect 8996 7828 9002 7880
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9456 7840 9505 7868
rect 9456 7828 9462 7840
rect 9493 7837 9505 7840
rect 9539 7837 9551 7871
rect 9493 7831 9551 7837
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7868 9643 7871
rect 9674 7868 9680 7880
rect 9631 7840 9680 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10042 7877 10048 7880
rect 10012 7871 10048 7877
rect 10012 7837 10024 7871
rect 10012 7831 10048 7837
rect 10042 7828 10048 7831
rect 10100 7828 10106 7880
rect 10134 7828 10140 7880
rect 10192 7868 10198 7880
rect 10229 7871 10287 7877
rect 10229 7868 10241 7871
rect 10192 7840 10241 7868
rect 10192 7828 10198 7840
rect 10229 7837 10241 7840
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 10962 7868 10968 7880
rect 10643 7840 10968 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 10962 7828 10968 7840
rect 11020 7828 11026 7880
rect 7374 7800 7380 7812
rect 7116 7772 7380 7800
rect 7009 7763 7067 7769
rect 7374 7760 7380 7772
rect 7432 7760 7438 7812
rect 7834 7760 7840 7812
rect 7892 7760 7898 7812
rect 3559 7704 4384 7732
rect 3559 7701 3571 7704
rect 3513 7695 3571 7701
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 4890 7732 4896 7744
rect 4672 7704 4896 7732
rect 4672 7692 4678 7704
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 7469 7735 7527 7741
rect 7469 7701 7481 7735
rect 7515 7732 7527 7735
rect 8404 7732 8432 7828
rect 9232 7800 9260 7828
rect 10321 7803 10379 7809
rect 10321 7800 10333 7803
rect 9232 7772 10333 7800
rect 10321 7769 10333 7772
rect 10367 7769 10379 7803
rect 11517 7803 11575 7809
rect 11517 7800 11529 7803
rect 10321 7763 10379 7769
rect 11164 7772 11529 7800
rect 7515 7704 8432 7732
rect 7515 7701 7527 7704
rect 7469 7695 7527 7701
rect 9030 7692 9036 7744
rect 9088 7692 9094 7744
rect 9953 7735 10011 7741
rect 9953 7701 9965 7735
rect 9999 7732 10011 7735
rect 10502 7732 10508 7744
rect 9999 7704 10508 7732
rect 9999 7701 10011 7704
rect 9953 7695 10011 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 11164 7741 11192 7772
rect 11517 7769 11529 7772
rect 11563 7769 11575 7803
rect 11517 7763 11575 7769
rect 12250 7760 12256 7812
rect 12308 7760 12314 7812
rect 13464 7800 13492 7899
rect 14366 7896 14372 7908
rect 14424 7936 14430 7948
rect 15856 7936 15884 8044
rect 18325 8041 18337 8044
rect 18371 8041 18383 8075
rect 18325 8035 18383 8041
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 17313 8007 17371 8013
rect 16632 7976 16712 8004
rect 16632 7964 16638 7976
rect 16684 7945 16712 7976
rect 17313 7973 17325 8007
rect 17359 8004 17371 8007
rect 17402 8004 17408 8016
rect 17359 7976 17408 8004
rect 17359 7973 17371 7976
rect 17313 7967 17371 7973
rect 17402 7964 17408 7976
rect 17460 7964 17466 8016
rect 17494 7964 17500 8016
rect 17552 7964 17558 8016
rect 14424 7908 15884 7936
rect 14424 7896 14430 7908
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 14826 7828 14832 7880
rect 14884 7868 14890 7880
rect 14921 7871 14979 7877
rect 14921 7868 14933 7871
rect 14884 7840 14933 7868
rect 14884 7828 14890 7840
rect 14921 7837 14933 7840
rect 14967 7837 14979 7871
rect 15562 7868 15568 7880
rect 14921 7831 14979 7837
rect 15028 7840 15568 7868
rect 14550 7800 14556 7812
rect 13464 7772 14556 7800
rect 14550 7760 14556 7772
rect 14608 7800 14614 7812
rect 15028 7800 15056 7840
rect 15562 7828 15568 7840
rect 15620 7828 15626 7880
rect 15749 7871 15807 7877
rect 15749 7837 15761 7871
rect 15795 7868 15807 7871
rect 15856 7868 15884 7908
rect 16669 7939 16727 7945
rect 16669 7905 16681 7939
rect 16715 7905 16727 7939
rect 16669 7899 16727 7905
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17862 7936 17868 7948
rect 17276 7908 17868 7936
rect 17276 7896 17282 7908
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 15795 7840 15884 7868
rect 15795 7837 15807 7840
rect 15749 7831 15807 7837
rect 16022 7828 16028 7880
rect 16080 7828 16086 7880
rect 16114 7828 16120 7880
rect 16172 7868 16178 7880
rect 16298 7868 16304 7880
rect 16172 7840 16304 7868
rect 16172 7828 16178 7840
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 14608 7772 15056 7800
rect 14608 7760 14614 7772
rect 15470 7760 15476 7812
rect 15528 7760 15534 7812
rect 15933 7803 15991 7809
rect 15933 7769 15945 7803
rect 15979 7800 15991 7803
rect 16408 7800 16436 7831
rect 16574 7828 16580 7880
rect 16632 7868 16638 7880
rect 16632 7840 17080 7868
rect 16632 7828 16638 7840
rect 17052 7800 17080 7840
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 17420 7800 17448 7831
rect 17494 7828 17500 7880
rect 17552 7868 17558 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17552 7840 18061 7868
rect 17552 7828 17558 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18414 7828 18420 7880
rect 18472 7828 18478 7880
rect 17681 7803 17739 7809
rect 17681 7800 17693 7803
rect 15979 7772 16436 7800
rect 16500 7772 16896 7800
rect 17052 7772 17693 7800
rect 15979 7769 15991 7772
rect 15933 7763 15991 7769
rect 10965 7735 11023 7741
rect 10965 7732 10977 7735
rect 10652 7704 10977 7732
rect 10652 7692 10658 7704
rect 10965 7701 10977 7704
rect 11011 7701 11023 7735
rect 10965 7695 11023 7701
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7701 11207 7735
rect 11149 7695 11207 7701
rect 12342 7692 12348 7744
rect 12400 7732 12406 7744
rect 12989 7735 13047 7741
rect 12989 7732 13001 7735
rect 12400 7704 13001 7732
rect 12400 7692 12406 7704
rect 12989 7701 13001 7704
rect 13035 7701 13047 7735
rect 12989 7695 13047 7701
rect 13262 7692 13268 7744
rect 13320 7692 13326 7744
rect 13446 7692 13452 7744
rect 13504 7732 13510 7744
rect 13722 7732 13728 7744
rect 13504 7704 13728 7732
rect 13504 7692 13510 7704
rect 13722 7692 13728 7704
rect 13780 7732 13786 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 13780 7704 13921 7732
rect 13780 7692 13786 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 14829 7735 14887 7741
rect 14829 7701 14841 7735
rect 14875 7732 14887 7735
rect 14918 7732 14924 7744
rect 14875 7704 14924 7732
rect 14875 7701 14887 7704
rect 14829 7695 14887 7701
rect 14918 7692 14924 7704
rect 14976 7732 14982 7744
rect 15948 7732 15976 7763
rect 14976 7704 15976 7732
rect 14976 7692 14982 7704
rect 16206 7692 16212 7744
rect 16264 7692 16270 7744
rect 16298 7692 16304 7744
rect 16356 7732 16362 7744
rect 16500 7732 16528 7772
rect 16356 7704 16528 7732
rect 16577 7735 16635 7741
rect 16356 7692 16362 7704
rect 16577 7701 16589 7735
rect 16623 7732 16635 7735
rect 16758 7732 16764 7744
rect 16623 7704 16764 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 16758 7692 16764 7704
rect 16816 7692 16822 7744
rect 16868 7732 16896 7772
rect 17681 7769 17693 7772
rect 17727 7769 17739 7803
rect 17681 7763 17739 7769
rect 17865 7803 17923 7809
rect 17865 7769 17877 7803
rect 17911 7769 17923 7803
rect 17865 7763 17923 7769
rect 17880 7732 17908 7763
rect 16868 7704 17908 7732
rect 1104 7642 18860 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 18860 7642
rect 1104 7568 18860 7590
rect 2869 7531 2927 7537
rect 2869 7497 2881 7531
rect 2915 7528 2927 7531
rect 3326 7528 3332 7540
rect 2915 7500 3332 7528
rect 2915 7497 2927 7500
rect 2869 7491 2927 7497
rect 3326 7488 3332 7500
rect 3384 7488 3390 7540
rect 5261 7531 5319 7537
rect 5261 7497 5273 7531
rect 5307 7528 5319 7531
rect 5810 7528 5816 7540
rect 5307 7500 5816 7528
rect 5307 7497 5319 7500
rect 5261 7491 5319 7497
rect 5810 7488 5816 7500
rect 5868 7488 5874 7540
rect 6641 7531 6699 7537
rect 6641 7497 6653 7531
rect 6687 7528 6699 7531
rect 6730 7528 6736 7540
rect 6687 7500 6736 7528
rect 6687 7497 6699 7500
rect 6641 7491 6699 7497
rect 6730 7488 6736 7500
rect 6788 7528 6794 7540
rect 9030 7528 9036 7540
rect 6788 7500 9036 7528
rect 6788 7488 6794 7500
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9398 7488 9404 7540
rect 9456 7488 9462 7540
rect 10870 7488 10876 7540
rect 10928 7488 10934 7540
rect 10962 7488 10968 7540
rect 11020 7528 11026 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 11020 7500 11621 7528
rect 11020 7488 11026 7500
rect 11609 7497 11621 7500
rect 11655 7497 11667 7531
rect 11609 7491 11667 7497
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 12308 7500 12357 7528
rect 12308 7488 12314 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 13446 7488 13452 7540
rect 13504 7488 13510 7540
rect 13909 7531 13967 7537
rect 13909 7497 13921 7531
rect 13955 7528 13967 7531
rect 13998 7528 14004 7540
rect 13955 7500 14004 7528
rect 13955 7497 13967 7500
rect 13909 7491 13967 7497
rect 13998 7488 14004 7500
rect 14056 7488 14062 7540
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 15160 7500 15516 7528
rect 15160 7488 15166 7500
rect 4246 7420 4252 7472
rect 4304 7460 4310 7472
rect 5534 7460 5540 7472
rect 4304 7432 5540 7460
rect 4304 7420 4310 7432
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 6880 7432 7052 7460
rect 6880 7420 6886 7432
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2556 7364 2605 7392
rect 2556 7352 2562 7364
rect 2593 7361 2605 7364
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 2682 7352 2688 7404
rect 2740 7392 2746 7404
rect 2740 7364 2912 7392
rect 2740 7352 2746 7364
rect 2884 7333 2912 7364
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 4893 7395 4951 7401
rect 4893 7392 4905 7395
rect 4856 7364 4905 7392
rect 4856 7352 4862 7364
rect 4893 7361 4905 7364
rect 4939 7361 4951 7395
rect 4893 7355 4951 7361
rect 5184 7364 6868 7392
rect 2869 7327 2927 7333
rect 2869 7293 2881 7327
rect 2915 7324 2927 7327
rect 5184 7324 5212 7364
rect 2915 7296 5212 7324
rect 2915 7293 2927 7296
rect 2869 7287 2927 7293
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 2685 7259 2743 7265
rect 2685 7256 2697 7259
rect 2648 7228 2697 7256
rect 2648 7216 2654 7228
rect 2685 7225 2697 7228
rect 2731 7225 2743 7259
rect 5718 7256 5724 7268
rect 2685 7219 2743 7225
rect 5276 7228 5724 7256
rect 4706 7148 4712 7200
rect 4764 7188 4770 7200
rect 5276 7197 5304 7228
rect 5718 7216 5724 7228
rect 5776 7216 5782 7268
rect 6840 7256 6868 7364
rect 6914 7352 6920 7404
rect 6972 7352 6978 7404
rect 7024 7401 7052 7432
rect 9582 7420 9588 7472
rect 9640 7420 9646 7472
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 12066 7460 12072 7472
rect 11931 7432 12072 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 12158 7420 12164 7472
rect 12216 7420 12222 7472
rect 13262 7420 13268 7472
rect 13320 7460 13326 7472
rect 14458 7460 14464 7472
rect 13320 7432 14136 7460
rect 13320 7420 13326 7432
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7392 9367 7395
rect 9398 7392 9404 7404
rect 9355 7364 9404 7392
rect 9355 7361 9367 7364
rect 9309 7355 9367 7361
rect 9398 7352 9404 7364
rect 9456 7352 9462 7404
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 11974 7352 11980 7404
rect 12032 7352 12038 7404
rect 12176 7392 12204 7420
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 12176 7364 12265 7392
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 13724 7395 13782 7401
rect 13724 7361 13736 7395
rect 13770 7361 13782 7395
rect 13724 7355 13782 7361
rect 6931 7324 6959 7352
rect 7650 7324 7656 7336
rect 6931 7296 7656 7324
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 12161 7327 12219 7333
rect 12161 7293 12173 7327
rect 12207 7324 12219 7327
rect 12342 7324 12348 7336
rect 12207 7296 12348 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 13739 7324 13767 7355
rect 13814 7352 13820 7404
rect 13872 7352 13878 7404
rect 14108 7401 14136 7432
rect 14292 7432 14464 7460
rect 14292 7401 14320 7432
rect 14458 7420 14464 7432
rect 14516 7460 14522 7472
rect 15289 7463 15347 7469
rect 15289 7460 15301 7463
rect 14516 7432 15301 7460
rect 14516 7420 14522 7432
rect 15289 7429 15301 7432
rect 15335 7429 15347 7463
rect 15289 7423 15347 7429
rect 14093 7395 14151 7401
rect 14093 7361 14105 7395
rect 14139 7361 14151 7395
rect 14093 7355 14151 7361
rect 14277 7395 14335 7401
rect 14277 7361 14289 7395
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 14366 7352 14372 7404
rect 14424 7352 14430 7404
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 14918 7352 14924 7404
rect 14976 7352 14982 7404
rect 15488 7401 15516 7500
rect 16132 7500 17632 7528
rect 16132 7401 16160 7500
rect 17604 7472 17632 7500
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 18012 7500 18337 7528
rect 18012 7488 18018 7500
rect 18325 7497 18337 7500
rect 18371 7497 18383 7531
rect 18325 7491 18383 7497
rect 17494 7420 17500 7472
rect 17552 7420 17558 7472
rect 17586 7420 17592 7472
rect 17644 7460 17650 7472
rect 18141 7463 18199 7469
rect 18141 7460 18153 7463
rect 17644 7432 18153 7460
rect 17644 7420 17650 7432
rect 18141 7429 18153 7432
rect 18187 7429 18199 7463
rect 18141 7423 18199 7429
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7361 15255 7395
rect 15197 7355 15255 7361
rect 15473 7395 15531 7401
rect 15473 7361 15485 7395
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 15212 7324 15240 7355
rect 15657 7327 15715 7333
rect 15657 7324 15669 7327
rect 13739 7296 15056 7324
rect 15212 7296 15669 7324
rect 7834 7256 7840 7268
rect 6840 7228 7840 7256
rect 7834 7216 7840 7228
rect 7892 7216 7898 7268
rect 11974 7216 11980 7268
rect 12032 7256 12038 7268
rect 13814 7256 13820 7268
rect 12032 7228 13820 7256
rect 12032 7216 12038 7228
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 14090 7216 14096 7268
rect 14148 7256 14154 7268
rect 14185 7259 14243 7265
rect 14185 7256 14197 7259
rect 14148 7228 14197 7256
rect 14148 7216 14154 7228
rect 14185 7225 14197 7228
rect 14231 7256 14243 7259
rect 14645 7259 14703 7265
rect 14645 7256 14657 7259
rect 14231 7228 14657 7256
rect 14231 7225 14243 7228
rect 14185 7219 14243 7225
rect 14645 7225 14657 7228
rect 14691 7225 14703 7259
rect 15028 7256 15056 7296
rect 15657 7293 15669 7296
rect 15703 7324 15715 7327
rect 16025 7327 16083 7333
rect 16025 7324 16037 7327
rect 15703 7296 16037 7324
rect 15703 7293 15715 7296
rect 15657 7287 15715 7293
rect 16025 7293 16037 7296
rect 16071 7293 16083 7327
rect 16500 7324 16528 7355
rect 16666 7352 16672 7404
rect 16724 7352 16730 7404
rect 16758 7352 16764 7404
rect 16816 7352 16822 7404
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 17957 7395 18015 7401
rect 17957 7392 17969 7395
rect 17184 7364 17969 7392
rect 17184 7352 17190 7364
rect 17957 7361 17969 7364
rect 18003 7361 18015 7395
rect 17957 7355 18015 7361
rect 18046 7324 18052 7336
rect 16500 7296 18052 7324
rect 16025 7287 16083 7293
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 15470 7256 15476 7268
rect 15028 7228 15476 7256
rect 14645 7219 14703 7225
rect 15470 7216 15476 7228
rect 15528 7216 15534 7268
rect 16114 7216 16120 7268
rect 16172 7256 16178 7268
rect 16301 7259 16359 7265
rect 16301 7256 16313 7259
rect 16172 7228 16313 7256
rect 16172 7216 16178 7228
rect 16301 7225 16313 7228
rect 16347 7256 16359 7259
rect 17126 7256 17132 7268
rect 16347 7228 17132 7256
rect 16347 7225 16359 7228
rect 16301 7219 16359 7225
rect 17126 7216 17132 7228
rect 17184 7216 17190 7268
rect 17218 7216 17224 7268
rect 17276 7256 17282 7268
rect 17865 7259 17923 7265
rect 17276 7228 17540 7256
rect 17276 7216 17282 7228
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4764 7160 5273 7188
rect 4764 7148 4770 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5261 7151 5319 7157
rect 5442 7148 5448 7200
rect 5500 7148 5506 7200
rect 12158 7148 12164 7200
rect 12216 7188 12222 7200
rect 12618 7188 12624 7200
rect 12216 7160 12624 7188
rect 12216 7148 12222 7160
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 13832 7188 13860 7216
rect 15010 7188 15016 7200
rect 13832 7160 15016 7188
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15102 7148 15108 7200
rect 15160 7148 15166 7200
rect 15378 7148 15384 7200
rect 15436 7188 15442 7200
rect 16945 7191 17003 7197
rect 16945 7188 16957 7191
rect 15436 7160 16957 7188
rect 15436 7148 15442 7160
rect 16945 7157 16957 7160
rect 16991 7157 17003 7191
rect 16945 7151 17003 7157
rect 17310 7148 17316 7200
rect 17368 7148 17374 7200
rect 17512 7197 17540 7228
rect 17865 7225 17877 7259
rect 17911 7256 17923 7259
rect 17954 7256 17960 7268
rect 17911 7228 17960 7256
rect 17911 7225 17923 7228
rect 17865 7219 17923 7225
rect 17954 7216 17960 7228
rect 18012 7216 18018 7268
rect 17497 7191 17555 7197
rect 17497 7157 17509 7191
rect 17543 7157 17555 7191
rect 17497 7151 17555 7157
rect 1104 7098 18860 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 18860 7098
rect 1104 7024 18860 7046
rect 5064 6987 5122 6993
rect 5064 6953 5076 6987
rect 5110 6984 5122 6987
rect 5442 6984 5448 6996
rect 5110 6956 5448 6984
rect 5110 6953 5122 6956
rect 5064 6947 5122 6953
rect 5442 6944 5448 6956
rect 5500 6944 5506 6996
rect 6178 6944 6184 6996
rect 6236 6984 6242 6996
rect 6549 6987 6607 6993
rect 6549 6984 6561 6987
rect 6236 6956 6561 6984
rect 6236 6944 6242 6956
rect 6549 6953 6561 6956
rect 6595 6953 6607 6987
rect 6549 6947 6607 6953
rect 11606 6944 11612 6996
rect 11664 6944 11670 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11992 6956 12081 6984
rect 9858 6876 9864 6928
rect 9916 6916 9922 6928
rect 11379 6919 11437 6925
rect 11379 6916 11391 6919
rect 9916 6888 11391 6916
rect 9916 6876 9922 6888
rect 11379 6885 11391 6888
rect 11425 6885 11437 6919
rect 11379 6879 11437 6885
rect 11517 6919 11575 6925
rect 11517 6885 11529 6919
rect 11563 6885 11575 6919
rect 11624 6916 11652 6944
rect 11992 6916 12020 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 12216 6956 12265 6984
rect 12216 6944 12222 6956
rect 12253 6953 12265 6956
rect 12299 6984 12311 6987
rect 12710 6984 12716 6996
rect 12299 6956 12716 6984
rect 12299 6953 12311 6956
rect 12253 6947 12311 6953
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 17037 6987 17095 6993
rect 17037 6953 17049 6987
rect 17083 6984 17095 6987
rect 17586 6984 17592 6996
rect 17083 6956 17592 6984
rect 17083 6953 17095 6956
rect 17037 6947 17095 6953
rect 11624 6888 12020 6916
rect 11517 6879 11575 6885
rect 4430 6808 4436 6860
rect 4488 6848 4494 6860
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 4488 6820 4813 6848
rect 4488 6808 4494 6820
rect 4801 6817 4813 6820
rect 4847 6848 4859 6851
rect 7098 6848 7104 6860
rect 4847 6820 7104 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 8570 6848 8576 6860
rect 8128 6820 8576 6848
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 6914 6780 6920 6792
rect 6871 6752 6920 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 6914 6740 6920 6752
rect 6972 6780 6978 6792
rect 8128 6780 8156 6820
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 10042 6848 10048 6860
rect 9324 6820 10048 6848
rect 6972 6752 8156 6780
rect 6972 6740 6978 6752
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 9324 6789 9352 6820
rect 10042 6808 10048 6820
rect 10100 6848 10106 6860
rect 11532 6848 11560 6879
rect 16758 6876 16764 6928
rect 16816 6916 16822 6928
rect 16945 6919 17003 6925
rect 16945 6916 16957 6919
rect 16816 6888 16957 6916
rect 16816 6876 16822 6888
rect 16945 6885 16957 6888
rect 16991 6885 17003 6919
rect 16945 6879 17003 6885
rect 10100 6820 10272 6848
rect 10100 6808 10106 6820
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 8260 6752 9321 6780
rect 8260 6740 8266 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 9858 6740 9864 6792
rect 9916 6740 9922 6792
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6749 10195 6783
rect 10137 6743 10195 6749
rect 4522 6672 4528 6724
rect 4580 6672 4586 6724
rect 4709 6715 4767 6721
rect 4709 6681 4721 6715
rect 4755 6712 4767 6715
rect 4798 6712 4804 6724
rect 4755 6684 4804 6712
rect 4755 6681 4767 6684
rect 4709 6675 4767 6681
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 6302 6684 6745 6712
rect 6733 6681 6745 6684
rect 6779 6681 6791 6715
rect 6733 6675 6791 6681
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 9582 6712 9588 6724
rect 8803 6684 9588 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 9582 6672 9588 6684
rect 9640 6672 9646 6724
rect 10152 6712 10180 6743
rect 9692 6684 10180 6712
rect 10244 6712 10272 6820
rect 10428 6820 11560 6848
rect 10428 6792 10456 6820
rect 11606 6808 11612 6860
rect 11664 6808 11670 6860
rect 16574 6848 16580 6860
rect 12176 6820 16580 6848
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10778 6740 10784 6792
rect 10836 6780 10842 6792
rect 12176 6790 12204 6820
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 11992 6789 12204 6790
rect 10873 6783 10931 6789
rect 10873 6780 10885 6783
rect 10836 6752 10885 6780
rect 10836 6740 10842 6752
rect 10873 6749 10885 6752
rect 10919 6749 10931 6783
rect 10873 6743 10931 6749
rect 11977 6783 12204 6789
rect 11977 6749 11989 6783
rect 12023 6762 12204 6783
rect 13165 6777 13223 6783
rect 13165 6774 13177 6777
rect 12023 6749 12035 6762
rect 11977 6743 12035 6749
rect 13096 6746 13177 6774
rect 11241 6715 11299 6721
rect 11241 6712 11253 6715
rect 10244 6684 11253 6712
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 4614 6644 4620 6656
rect 4387 6616 4620 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 9493 6647 9551 6653
rect 9493 6613 9505 6647
rect 9539 6644 9551 6647
rect 9692 6644 9720 6684
rect 11241 6681 11253 6684
rect 11287 6681 11299 6715
rect 11241 6675 11299 6681
rect 12066 6672 12072 6724
rect 12124 6712 12130 6724
rect 12437 6715 12495 6721
rect 12437 6712 12449 6715
rect 12124 6684 12449 6712
rect 12124 6672 12130 6684
rect 12437 6681 12449 6684
rect 12483 6681 12495 6715
rect 12437 6675 12495 6681
rect 9539 6616 9720 6644
rect 9539 6613 9551 6616
rect 9493 6607 9551 6613
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10410 6644 10416 6656
rect 9824 6616 10416 6644
rect 9824 6604 9830 6616
rect 10410 6604 10416 6616
rect 10468 6604 10474 6656
rect 11057 6647 11115 6653
rect 11057 6613 11069 6647
rect 11103 6644 11115 6647
rect 11146 6644 11152 6656
rect 11103 6616 11152 6644
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11146 6604 11152 6616
rect 11204 6604 11210 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12227 6647 12285 6653
rect 12227 6644 12239 6647
rect 11848 6616 12239 6644
rect 11848 6604 11854 6616
rect 12227 6613 12239 6616
rect 12273 6644 12285 6647
rect 12342 6644 12348 6656
rect 12273 6616 12348 6644
rect 12273 6613 12285 6616
rect 12227 6607 12285 6613
rect 12342 6604 12348 6616
rect 12400 6604 12406 6656
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 13096 6644 13124 6746
rect 13165 6743 13177 6746
rect 13211 6743 13223 6777
rect 13165 6737 13223 6743
rect 16666 6740 16672 6792
rect 16724 6740 16730 6792
rect 17052 6780 17080 6947
rect 17586 6944 17592 6956
rect 17644 6944 17650 6996
rect 16776 6752 17080 6780
rect 16776 6721 16804 6752
rect 17218 6740 17224 6792
rect 17276 6740 17282 6792
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 17681 6783 17739 6789
rect 17681 6780 17693 6783
rect 17368 6752 17693 6780
rect 17368 6740 17374 6752
rect 17681 6749 17693 6752
rect 17727 6749 17739 6783
rect 17681 6743 17739 6749
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6780 18199 6783
rect 18414 6780 18420 6792
rect 18187 6752 18420 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 16761 6715 16819 6721
rect 16761 6681 16773 6715
rect 16807 6681 16819 6715
rect 16761 6675 16819 6681
rect 16945 6715 17003 6721
rect 16945 6681 16957 6715
rect 16991 6712 17003 6715
rect 17328 6712 17356 6740
rect 16991 6684 17356 6712
rect 16991 6681 17003 6684
rect 16945 6675 17003 6681
rect 12676 6616 13124 6644
rect 13265 6647 13323 6653
rect 12676 6604 12682 6616
rect 13265 6613 13277 6647
rect 13311 6644 13323 6647
rect 13446 6644 13452 6656
rect 13311 6616 13452 6644
rect 13311 6613 13323 6616
rect 13265 6607 13323 6613
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 15010 6604 15016 6656
rect 15068 6644 15074 6656
rect 16206 6644 16212 6656
rect 15068 6616 16212 6644
rect 15068 6604 15074 6616
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 17310 6604 17316 6656
rect 17368 6604 17374 6656
rect 1104 6554 18860 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 18860 6554
rect 1104 6480 18860 6502
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 6181 6443 6239 6449
rect 6181 6440 6193 6443
rect 4580 6412 6193 6440
rect 4580 6400 4586 6412
rect 6181 6409 6193 6412
rect 6227 6409 6239 6443
rect 6914 6440 6920 6452
rect 6181 6403 6239 6409
rect 6564 6412 6920 6440
rect 6457 6375 6515 6381
rect 6457 6372 6469 6375
rect 5934 6344 6469 6372
rect 6457 6341 6469 6344
rect 6503 6341 6515 6375
rect 6457 6335 6515 6341
rect 4430 6264 4436 6316
rect 4488 6264 4494 6316
rect 6564 6313 6592 6412
rect 6914 6400 6920 6412
rect 6972 6400 6978 6452
rect 7561 6443 7619 6449
rect 7561 6409 7573 6443
rect 7607 6440 7619 6443
rect 8110 6440 8116 6452
rect 7607 6412 8116 6440
rect 7607 6409 7619 6412
rect 7561 6403 7619 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 8812 6412 9260 6440
rect 8812 6400 8818 6412
rect 7101 6375 7159 6381
rect 7101 6372 7113 6375
rect 6748 6344 7113 6372
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 4709 6239 4767 6245
rect 4709 6205 4721 6239
rect 4755 6236 4767 6239
rect 4798 6236 4804 6248
rect 4755 6208 4804 6236
rect 4755 6205 4767 6208
rect 4709 6199 4767 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 2958 6060 2964 6112
rect 3016 6100 3022 6112
rect 6748 6100 6776 6344
rect 7101 6341 7113 6344
rect 7147 6341 7159 6375
rect 7101 6335 7159 6341
rect 7926 6332 7932 6384
rect 7984 6372 7990 6384
rect 9232 6381 9260 6412
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 10505 6443 10563 6449
rect 10505 6440 10517 6443
rect 9364 6412 10517 6440
rect 9364 6400 9370 6412
rect 10505 6409 10517 6412
rect 10551 6409 10563 6443
rect 10505 6403 10563 6409
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 11606 6440 11612 6452
rect 10836 6412 11612 6440
rect 10836 6400 10842 6412
rect 11606 6400 11612 6412
rect 11664 6400 11670 6452
rect 12069 6443 12127 6449
rect 12069 6409 12081 6443
rect 12115 6440 12127 6443
rect 12115 6412 12480 6440
rect 12115 6409 12127 6412
rect 12069 6403 12127 6409
rect 9217 6375 9275 6381
rect 7984 6344 8433 6372
rect 7984 6332 7990 6344
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6304 7343 6307
rect 7650 6304 7656 6316
rect 7331 6276 7656 6304
rect 7331 6273 7343 6276
rect 7285 6267 7343 6273
rect 7650 6264 7656 6276
rect 7708 6264 7714 6316
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6304 7803 6307
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 7791 6276 8217 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7760 6236 7788 6267
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8405 6304 8433 6344
rect 9217 6341 9229 6375
rect 9263 6372 9275 6375
rect 9950 6372 9956 6384
rect 9263 6344 9956 6372
rect 9263 6341 9275 6344
rect 9217 6335 9275 6341
rect 9950 6332 9956 6344
rect 10008 6332 10014 6384
rect 10321 6375 10379 6381
rect 10321 6341 10333 6375
rect 10367 6372 10379 6375
rect 11885 6375 11943 6381
rect 10367 6344 11008 6372
rect 10367 6341 10379 6344
rect 10321 6335 10379 6341
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8405 6302 8524 6304
rect 8570 6302 8585 6304
rect 8405 6276 8585 6302
rect 8496 6274 8585 6276
rect 8573 6273 8585 6274
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6304 8723 6307
rect 8711 6276 8800 6304
rect 8711 6273 8723 6276
rect 8665 6267 8723 6273
rect 6963 6208 7788 6236
rect 7929 6239 7987 6245
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8312 6236 8340 6264
rect 7975 6208 8340 6236
rect 8772 6236 8800 6276
rect 8846 6264 8852 6316
rect 8904 6264 8910 6316
rect 8938 6264 8944 6316
rect 8996 6304 9002 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8996 6276 9137 6304
rect 8996 6264 9002 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 9125 6267 9183 6273
rect 9766 6264 9772 6316
rect 9824 6304 9830 6316
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 9824 6276 9873 6304
rect 9824 6264 9830 6276
rect 9861 6273 9873 6276
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 10042 6264 10048 6316
rect 10100 6264 10106 6316
rect 10137 6307 10195 6313
rect 10137 6273 10149 6307
rect 10183 6273 10195 6307
rect 10137 6267 10195 6273
rect 9033 6239 9091 6245
rect 8772 6208 8892 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8864 6180 8892 6208
rect 9033 6205 9045 6239
rect 9079 6236 9091 6239
rect 10152 6236 10180 6267
rect 10226 6264 10232 6316
rect 10284 6304 10290 6316
rect 10413 6307 10471 6313
rect 10413 6304 10425 6307
rect 10284 6276 10425 6304
rect 10284 6264 10290 6276
rect 10413 6273 10425 6276
rect 10459 6273 10471 6307
rect 10413 6267 10471 6273
rect 10686 6264 10692 6316
rect 10744 6264 10750 6316
rect 10980 6313 11008 6344
rect 11885 6341 11897 6375
rect 11931 6372 11943 6375
rect 11974 6372 11980 6384
rect 11931 6344 11980 6372
rect 11931 6341 11943 6344
rect 11885 6335 11943 6341
rect 11974 6332 11980 6344
rect 12032 6332 12038 6384
rect 12452 6381 12480 6412
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 13909 6443 13967 6449
rect 13909 6440 13921 6443
rect 13872 6412 13921 6440
rect 13872 6400 13878 6412
rect 13909 6409 13921 6412
rect 13955 6409 13967 6443
rect 13909 6403 13967 6409
rect 15930 6400 15936 6452
rect 15988 6440 15994 6452
rect 16393 6443 16451 6449
rect 16393 6440 16405 6443
rect 15988 6412 16405 6440
rect 15988 6400 15994 6412
rect 16393 6409 16405 6412
rect 16439 6409 16451 6443
rect 16393 6403 16451 6409
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6409 17095 6443
rect 17037 6403 17095 6409
rect 12437 6375 12495 6381
rect 12437 6341 12449 6375
rect 12483 6341 12495 6375
rect 12437 6335 12495 6341
rect 13446 6332 13452 6384
rect 13504 6332 13510 6384
rect 15197 6375 15255 6381
rect 15197 6341 15209 6375
rect 15243 6372 15255 6375
rect 15470 6372 15476 6384
rect 15243 6344 15476 6372
rect 15243 6341 15255 6344
rect 15197 6335 15255 6341
rect 15470 6332 15476 6344
rect 15528 6372 15534 6384
rect 17052 6372 17080 6403
rect 15528 6344 17080 6372
rect 15528 6332 15534 6344
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11514 6264 11520 6316
rect 11572 6264 11578 6316
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 15013 6307 15071 6313
rect 15013 6304 15025 6307
rect 14884 6276 15025 6304
rect 14884 6264 14890 6276
rect 15013 6273 15025 6276
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 10778 6236 10784 6248
rect 9079 6208 9904 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 9876 6180 9904 6208
rect 10060 6208 10784 6236
rect 10060 6180 10088 6208
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 10870 6196 10876 6248
rect 10928 6236 10934 6248
rect 12161 6239 12219 6245
rect 12161 6236 12173 6239
rect 10928 6208 12173 6236
rect 10928 6196 10934 6208
rect 12161 6205 12173 6208
rect 12207 6236 12219 6239
rect 12526 6236 12532 6248
rect 12207 6208 12532 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 14550 6196 14556 6248
rect 14608 6236 14614 6248
rect 15102 6236 15108 6248
rect 14608 6208 15108 6236
rect 14608 6196 14614 6208
rect 15102 6196 15108 6208
rect 15160 6236 15166 6248
rect 15304 6236 15332 6267
rect 15378 6264 15384 6316
rect 15436 6264 15442 6316
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 15160 6208 15332 6236
rect 15160 6196 15166 6208
rect 15562 6196 15568 6248
rect 15620 6236 15626 6248
rect 15948 6236 15976 6267
rect 16206 6264 16212 6316
rect 16264 6264 16270 6316
rect 16298 6264 16304 6316
rect 16356 6264 16362 6316
rect 16482 6264 16488 6316
rect 16540 6264 16546 6316
rect 17402 6264 17408 6316
rect 17460 6304 17466 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 17460 6276 18245 6304
rect 17460 6264 17466 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 16390 6236 16396 6248
rect 15620 6208 16396 6236
rect 15620 6196 15626 6208
rect 16390 6196 16396 6208
rect 16448 6236 16454 6248
rect 16574 6236 16580 6248
rect 16448 6208 16580 6236
rect 16448 6196 16454 6208
rect 16574 6196 16580 6208
rect 16632 6196 16638 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 17276 6208 17325 6236
rect 17276 6196 17282 6208
rect 17313 6205 17325 6208
rect 17359 6236 17371 6239
rect 17494 6236 17500 6248
rect 17359 6208 17500 6236
rect 17359 6205 17371 6208
rect 17313 6199 17371 6205
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 18506 6196 18512 6248
rect 18564 6196 18570 6248
rect 8018 6128 8024 6180
rect 8076 6128 8082 6180
rect 8846 6128 8852 6180
rect 8904 6128 8910 6180
rect 9858 6128 9864 6180
rect 9916 6168 9922 6180
rect 9953 6171 10011 6177
rect 9953 6168 9965 6171
rect 9916 6140 9965 6168
rect 9916 6128 9922 6140
rect 9953 6137 9965 6140
rect 9999 6137 10011 6171
rect 9953 6131 10011 6137
rect 10042 6128 10048 6180
rect 10100 6128 10106 6180
rect 10594 6128 10600 6180
rect 10652 6168 10658 6180
rect 10652 6140 11928 6168
rect 10652 6128 10658 6140
rect 7282 6100 7288 6112
rect 3016 6072 7288 6100
rect 3016 6060 3022 6072
rect 7282 6060 7288 6072
rect 7340 6060 7346 6112
rect 7466 6060 7472 6112
rect 7524 6060 7530 6112
rect 8481 6103 8539 6109
rect 8481 6069 8493 6103
rect 8527 6100 8539 6103
rect 8662 6100 8668 6112
rect 8527 6072 8668 6100
rect 8527 6069 8539 6072
rect 8481 6063 8539 6069
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 10134 6100 10140 6112
rect 8812 6072 10140 6100
rect 8812 6060 8818 6072
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10502 6060 10508 6112
rect 10560 6100 10566 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10560 6072 10885 6100
rect 10560 6060 10566 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 10962 6060 10968 6112
rect 11020 6060 11026 6112
rect 11900 6109 11928 6140
rect 16022 6128 16028 6180
rect 16080 6168 16086 6180
rect 16117 6171 16175 6177
rect 16117 6168 16129 6171
rect 16080 6140 16129 6168
rect 16080 6128 16086 6140
rect 16117 6137 16129 6140
rect 16163 6168 16175 6171
rect 16163 6140 17356 6168
rect 16163 6137 16175 6140
rect 16117 6131 16175 6137
rect 17328 6112 17356 6140
rect 11885 6103 11943 6109
rect 11885 6069 11897 6103
rect 11931 6069 11943 6103
rect 11885 6063 11943 6069
rect 15562 6060 15568 6112
rect 15620 6060 15626 6112
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 15746 6100 15752 6112
rect 15703 6072 15752 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 15838 6060 15844 6112
rect 15896 6100 15902 6112
rect 16758 6100 16764 6112
rect 15896 6072 16764 6100
rect 15896 6060 15902 6072
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 17310 6060 17316 6112
rect 17368 6060 17374 6112
rect 1104 6010 18860 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 18860 6010
rect 1104 5936 18860 5958
rect 4706 5856 4712 5908
rect 4764 5856 4770 5908
rect 5258 5856 5264 5908
rect 5316 5896 5322 5908
rect 9122 5896 9128 5908
rect 5316 5868 9128 5896
rect 5316 5856 5322 5868
rect 9122 5856 9128 5868
rect 9180 5856 9186 5908
rect 9858 5896 9864 5908
rect 9232 5868 9864 5896
rect 4525 5831 4583 5837
rect 4525 5797 4537 5831
rect 4571 5828 4583 5831
rect 4798 5828 4804 5840
rect 4571 5800 4804 5828
rect 4571 5797 4583 5800
rect 4525 5791 4583 5797
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 5077 5831 5135 5837
rect 5077 5797 5089 5831
rect 5123 5828 5135 5831
rect 5350 5828 5356 5840
rect 5123 5800 5356 5828
rect 5123 5797 5135 5800
rect 5077 5791 5135 5797
rect 5350 5788 5356 5800
rect 5408 5788 5414 5840
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 7524 5800 7696 5828
rect 7524 5788 7530 5800
rect 7668 5769 7696 5800
rect 7742 5788 7748 5840
rect 7800 5828 7806 5840
rect 8389 5831 8447 5837
rect 7800 5800 8064 5828
rect 7800 5788 7806 5800
rect 7653 5763 7711 5769
rect 7653 5729 7665 5763
rect 7699 5760 7711 5763
rect 8036 5760 8064 5800
rect 8389 5797 8401 5831
rect 8435 5828 8447 5831
rect 9030 5828 9036 5840
rect 8435 5800 9036 5828
rect 8435 5797 8447 5800
rect 8389 5791 8447 5797
rect 9030 5788 9036 5800
rect 9088 5788 9094 5840
rect 8846 5760 8852 5772
rect 7699 5732 7972 5760
rect 8036 5732 8852 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 7282 5652 7288 5704
rect 7340 5652 7346 5704
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 7742 5692 7748 5704
rect 7515 5664 7748 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7944 5692 7972 5732
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7944 5664 8125 5692
rect 7837 5655 7895 5661
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 4709 5627 4767 5633
rect 4709 5593 4721 5627
rect 4755 5624 4767 5627
rect 4890 5624 4896 5636
rect 4755 5596 4896 5624
rect 4755 5593 4767 5596
rect 4709 5587 4767 5593
rect 4890 5584 4896 5596
rect 4948 5584 4954 5636
rect 7300 5556 7328 5652
rect 7377 5627 7435 5633
rect 7377 5593 7389 5627
rect 7423 5624 7435 5627
rect 7852 5624 7880 5655
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8260 5664 8493 5692
rect 8260 5652 8266 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 9232 5692 9260 5868
rect 9858 5856 9864 5868
rect 9916 5856 9922 5908
rect 10321 5899 10379 5905
rect 10321 5865 10333 5899
rect 10367 5896 10379 5899
rect 10962 5896 10968 5908
rect 10367 5868 10968 5896
rect 10367 5865 10379 5868
rect 10321 5859 10379 5865
rect 10134 5828 10140 5840
rect 9692 5800 10140 5828
rect 9692 5769 9720 5800
rect 10134 5788 10140 5800
rect 10192 5828 10198 5840
rect 10336 5828 10364 5859
rect 10962 5856 10968 5868
rect 11020 5856 11026 5908
rect 11974 5856 11980 5908
rect 12032 5856 12038 5908
rect 15105 5899 15163 5905
rect 15105 5865 15117 5899
rect 15151 5896 15163 5899
rect 15194 5896 15200 5908
rect 15151 5868 15200 5896
rect 15151 5865 15163 5868
rect 15105 5859 15163 5865
rect 15194 5856 15200 5868
rect 15252 5856 15258 5908
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5896 15347 5899
rect 15562 5896 15568 5908
rect 15335 5868 15568 5896
rect 15335 5865 15347 5868
rect 15289 5859 15347 5865
rect 15562 5856 15568 5868
rect 15620 5856 15626 5908
rect 16206 5856 16212 5908
rect 16264 5896 16270 5908
rect 16264 5868 16521 5896
rect 16264 5856 16270 5868
rect 10192 5800 10364 5828
rect 11149 5831 11207 5837
rect 10192 5788 10198 5800
rect 11149 5797 11161 5831
rect 11195 5828 11207 5831
rect 15381 5831 15439 5837
rect 11195 5800 15332 5828
rect 11195 5797 11207 5800
rect 11149 5791 11207 5797
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 9677 5723 9735 5729
rect 10045 5763 10103 5769
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10091 5732 10456 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 8711 5664 9260 5692
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 9585 5695 9643 5701
rect 9585 5661 9597 5695
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 9861 5695 9919 5701
rect 9861 5661 9873 5695
rect 9907 5692 9919 5695
rect 9950 5692 9956 5704
rect 9907 5664 9956 5692
rect 9907 5661 9919 5664
rect 9861 5655 9919 5661
rect 7423 5596 7880 5624
rect 8021 5627 8079 5633
rect 7423 5593 7435 5596
rect 7377 5587 7435 5593
rect 8021 5593 8033 5627
rect 8067 5624 8079 5627
rect 8294 5624 8300 5636
rect 8067 5596 8300 5624
rect 8067 5593 8079 5596
rect 8021 5587 8079 5593
rect 8294 5584 8300 5596
rect 8352 5584 8358 5636
rect 8386 5584 8392 5636
rect 8444 5624 8450 5636
rect 8573 5627 8631 5633
rect 8573 5624 8585 5627
rect 8444 5596 8585 5624
rect 8444 5584 8450 5596
rect 8573 5593 8585 5596
rect 8619 5593 8631 5627
rect 8573 5587 8631 5593
rect 8754 5584 8760 5636
rect 8812 5624 8818 5636
rect 9600 5624 9628 5655
rect 9950 5652 9956 5664
rect 10008 5692 10014 5704
rect 10229 5695 10287 5701
rect 10229 5692 10241 5695
rect 10008 5664 10241 5692
rect 10008 5652 10014 5664
rect 10229 5661 10241 5664
rect 10275 5692 10287 5695
rect 10318 5692 10324 5704
rect 10275 5664 10324 5692
rect 10275 5661 10287 5664
rect 10229 5655 10287 5661
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 8812 5596 9628 5624
rect 8812 5584 8818 5596
rect 9674 5584 9680 5636
rect 9732 5624 9738 5636
rect 10042 5624 10048 5636
rect 9732 5596 10048 5624
rect 9732 5584 9738 5596
rect 10042 5584 10048 5596
rect 10100 5584 10106 5636
rect 10428 5624 10456 5732
rect 10870 5720 10876 5772
rect 10928 5760 10934 5772
rect 10965 5763 11023 5769
rect 10965 5760 10977 5763
rect 10928 5732 10977 5760
rect 10928 5720 10934 5732
rect 10965 5729 10977 5732
rect 11011 5729 11023 5763
rect 10965 5723 11023 5729
rect 12342 5720 12348 5772
rect 12400 5760 12406 5772
rect 14645 5763 14703 5769
rect 12400 5732 14136 5760
rect 12400 5720 12406 5732
rect 10502 5652 10508 5704
rect 10560 5652 10566 5704
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 10612 5664 10793 5692
rect 10612 5624 10640 5664
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 11149 5695 11207 5701
rect 11149 5661 11161 5695
rect 11195 5661 11207 5695
rect 11149 5655 11207 5661
rect 10428 5596 10640 5624
rect 10689 5627 10747 5633
rect 10689 5593 10701 5627
rect 10735 5624 10747 5627
rect 11164 5624 11192 5655
rect 12066 5652 12072 5704
rect 12124 5692 12130 5704
rect 12636 5701 12664 5732
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 12124 5664 12173 5692
rect 12124 5652 12130 5664
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 12768 5664 13492 5692
rect 12768 5652 12774 5664
rect 10735 5596 11192 5624
rect 10735 5593 10747 5596
rect 10689 5587 10747 5593
rect 12250 5584 12256 5636
rect 12308 5624 12314 5636
rect 12345 5627 12403 5633
rect 12345 5624 12357 5627
rect 12308 5596 12357 5624
rect 12308 5584 12314 5596
rect 12345 5593 12357 5596
rect 12391 5624 12403 5627
rect 12437 5627 12495 5633
rect 12437 5624 12449 5627
rect 12391 5596 12449 5624
rect 12391 5593 12403 5596
rect 12345 5587 12403 5593
rect 12437 5593 12449 5596
rect 12483 5593 12495 5627
rect 12437 5587 12495 5593
rect 12989 5627 13047 5633
rect 12989 5593 13001 5627
rect 13035 5593 13047 5627
rect 13464 5624 13492 5664
rect 13538 5652 13544 5704
rect 13596 5652 13602 5704
rect 14108 5701 14136 5732
rect 14645 5729 14657 5763
rect 14691 5760 14703 5763
rect 15194 5760 15200 5772
rect 14691 5732 15200 5760
rect 14691 5729 14703 5732
rect 14645 5723 14703 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 15304 5760 15332 5800
rect 15381 5797 15393 5831
rect 15427 5828 15439 5831
rect 15841 5831 15899 5837
rect 15841 5828 15853 5831
rect 15427 5800 15853 5828
rect 15427 5797 15439 5800
rect 15381 5791 15439 5797
rect 15841 5797 15853 5800
rect 15887 5797 15899 5831
rect 15841 5791 15899 5797
rect 16390 5788 16396 5840
rect 16448 5788 16454 5840
rect 15654 5760 15660 5772
rect 15304 5732 15660 5760
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15746 5720 15752 5772
rect 15804 5720 15810 5772
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15378 5692 15384 5704
rect 14783 5664 15384 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15930 5652 15936 5704
rect 15988 5701 15994 5704
rect 15988 5695 16037 5701
rect 15988 5661 15991 5695
rect 16025 5661 16037 5695
rect 15988 5655 16037 5661
rect 15988 5652 15994 5655
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 16408 5701 16436 5788
rect 16493 5701 16521 5868
rect 17034 5856 17040 5908
rect 17092 5896 17098 5908
rect 18325 5899 18383 5905
rect 18325 5896 18337 5899
rect 17092 5868 18337 5896
rect 17092 5856 17098 5868
rect 18325 5865 18337 5868
rect 18371 5865 18383 5899
rect 18325 5859 18383 5865
rect 16392 5695 16450 5701
rect 16172 5664 16217 5692
rect 16172 5652 16178 5664
rect 16392 5661 16404 5695
rect 16438 5661 16450 5695
rect 16392 5655 16450 5661
rect 16478 5695 16536 5701
rect 16478 5661 16490 5695
rect 16524 5661 16536 5695
rect 16478 5655 16536 5661
rect 16574 5652 16580 5704
rect 16632 5652 16638 5704
rect 16758 5652 16764 5704
rect 16816 5652 16822 5704
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5692 17003 5695
rect 17310 5692 17316 5704
rect 16991 5664 17316 5692
rect 16991 5661 17003 5664
rect 16945 5655 17003 5661
rect 17310 5652 17316 5664
rect 17368 5652 17374 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 18598 5692 18604 5704
rect 18555 5664 18604 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 14277 5627 14335 5633
rect 14277 5624 14289 5627
rect 13464 5596 14289 5624
rect 12989 5587 13047 5593
rect 14277 5593 14289 5596
rect 14323 5624 14335 5627
rect 14642 5624 14648 5636
rect 14323 5596 14648 5624
rect 14323 5593 14335 5596
rect 14277 5587 14335 5593
rect 8110 5556 8116 5568
rect 7300 5528 8116 5556
rect 8110 5516 8116 5528
rect 8168 5516 8174 5568
rect 8205 5559 8263 5565
rect 8205 5525 8217 5559
rect 8251 5556 8263 5559
rect 8478 5556 8484 5568
rect 8251 5528 8484 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 8478 5516 8484 5528
rect 8536 5556 8542 5568
rect 8662 5556 8668 5568
rect 8536 5528 8668 5556
rect 8536 5516 8542 5528
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 10778 5556 10784 5568
rect 9180 5528 10784 5556
rect 9180 5516 9186 5528
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 10870 5516 10876 5568
rect 10928 5516 10934 5568
rect 12158 5516 12164 5568
rect 12216 5556 12222 5568
rect 13004 5556 13032 5587
rect 14642 5584 14648 5596
rect 14700 5584 14706 5636
rect 16209 5627 16267 5633
rect 16209 5593 16221 5627
rect 16255 5624 16267 5627
rect 16776 5624 16804 5652
rect 16255 5596 16380 5624
rect 16255 5593 16267 5596
rect 16209 5587 16267 5593
rect 12216 5528 13032 5556
rect 12216 5516 12222 5528
rect 14458 5516 14464 5568
rect 14516 5516 14522 5568
rect 16352 5556 16380 5596
rect 16500 5596 16804 5624
rect 16500 5556 16528 5596
rect 16850 5584 16856 5636
rect 16908 5584 16914 5636
rect 16352 5528 16528 5556
rect 17126 5516 17132 5568
rect 17184 5516 17190 5568
rect 1104 5466 18860 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 18860 5466
rect 1104 5392 18860 5414
rect 9217 5355 9275 5361
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 10226 5352 10232 5364
rect 9263 5324 10232 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 10226 5312 10232 5324
rect 10284 5352 10290 5364
rect 10413 5355 10471 5361
rect 10284 5324 10364 5352
rect 10284 5312 10290 5324
rect 4801 5287 4859 5293
rect 4801 5253 4813 5287
rect 4847 5284 4859 5287
rect 5534 5284 5540 5296
rect 4847 5256 5540 5284
rect 4847 5253 4859 5256
rect 4801 5247 4859 5253
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5216 5043 5219
rect 5261 5219 5319 5225
rect 5261 5216 5273 5219
rect 5031 5188 5273 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5261 5185 5273 5188
rect 5307 5216 5319 5219
rect 5350 5216 5356 5228
rect 5307 5188 5356 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 5460 5225 5488 5256
rect 5534 5244 5540 5256
rect 5592 5244 5598 5296
rect 8294 5244 8300 5296
rect 8352 5284 8358 5296
rect 8849 5287 8907 5293
rect 8849 5284 8861 5287
rect 8352 5256 8861 5284
rect 8352 5244 8358 5256
rect 8849 5253 8861 5256
rect 8895 5284 8907 5287
rect 9490 5284 9496 5296
rect 8895 5256 9496 5284
rect 8895 5253 8907 5256
rect 8849 5247 8907 5253
rect 9490 5244 9496 5256
rect 9548 5244 9554 5296
rect 9950 5244 9956 5296
rect 10008 5244 10014 5296
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5216 5503 5219
rect 5491 5188 5525 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 7926 5176 7932 5228
rect 7984 5216 7990 5228
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 7984 5188 8217 5216
rect 7984 5176 7990 5188
rect 8205 5185 8217 5188
rect 8251 5216 8263 5219
rect 8478 5216 8484 5228
rect 8251 5188 8484 5216
rect 8251 5185 8263 5188
rect 8205 5179 8263 5185
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5216 8723 5219
rect 8754 5216 8760 5228
rect 8711 5188 8760 5216
rect 8711 5185 8723 5188
rect 8665 5179 8723 5185
rect 8754 5176 8760 5188
rect 8812 5176 8818 5228
rect 8938 5176 8944 5228
rect 8996 5176 9002 5228
rect 9030 5176 9036 5228
rect 9088 5176 9094 5228
rect 9398 5176 9404 5228
rect 9456 5216 9462 5228
rect 9677 5219 9735 5225
rect 9677 5216 9689 5219
rect 9456 5188 9689 5216
rect 9456 5176 9462 5188
rect 9677 5185 9689 5188
rect 9723 5185 9735 5219
rect 9677 5179 9735 5185
rect 9861 5219 9919 5225
rect 9861 5185 9873 5219
rect 9907 5185 9919 5219
rect 9861 5179 9919 5185
rect 10045 5219 10103 5225
rect 10045 5185 10057 5219
rect 10091 5216 10103 5219
rect 10134 5216 10140 5228
rect 10091 5188 10140 5216
rect 10091 5185 10103 5188
rect 10045 5179 10103 5185
rect 8113 5151 8171 5157
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 8386 5148 8392 5160
rect 8159 5120 8392 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8496 5148 8524 5176
rect 9582 5148 9588 5160
rect 8496 5120 9588 5148
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 8573 5083 8631 5089
rect 8573 5049 8585 5083
rect 8619 5080 8631 5083
rect 9030 5080 9036 5092
rect 8619 5052 9036 5080
rect 8619 5049 8631 5052
rect 8573 5043 8631 5049
rect 9030 5040 9036 5052
rect 9088 5080 9094 5092
rect 9876 5080 9904 5179
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10336 5225 10364 5324
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 10870 5352 10876 5364
rect 10459 5324 10876 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 10870 5312 10876 5324
rect 10928 5312 10934 5364
rect 15565 5355 15623 5361
rect 15565 5321 15577 5355
rect 15611 5352 15623 5355
rect 15746 5352 15752 5364
rect 15611 5324 15752 5352
rect 15611 5321 15623 5324
rect 15565 5315 15623 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16114 5312 16120 5364
rect 16172 5312 16178 5364
rect 16301 5355 16359 5361
rect 16301 5321 16313 5355
rect 16347 5352 16359 5355
rect 16482 5352 16488 5364
rect 16347 5324 16488 5352
rect 16347 5321 16359 5324
rect 16301 5315 16359 5321
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 12158 5244 12164 5296
rect 12216 5284 12222 5296
rect 12345 5287 12403 5293
rect 12345 5284 12357 5287
rect 12216 5256 12357 5284
rect 12216 5244 12222 5256
rect 12345 5253 12357 5256
rect 12391 5253 12403 5287
rect 12345 5247 12403 5253
rect 13630 5244 13636 5296
rect 13688 5244 13694 5296
rect 14642 5244 14648 5296
rect 14700 5244 14706 5296
rect 15470 5284 15476 5296
rect 15028 5256 15476 5284
rect 10321 5219 10379 5225
rect 10321 5185 10333 5219
rect 10367 5185 10379 5219
rect 10321 5179 10379 5185
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5216 10563 5219
rect 10686 5216 10692 5228
rect 10551 5188 10692 5216
rect 10551 5185 10563 5188
rect 10505 5179 10563 5185
rect 9088 5052 9904 5080
rect 10229 5083 10287 5089
rect 9088 5040 9094 5052
rect 10229 5049 10241 5083
rect 10275 5080 10287 5083
rect 10520 5080 10548 5179
rect 10686 5176 10692 5188
rect 10744 5176 10750 5228
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12250 5216 12256 5228
rect 12023 5188 12256 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12250 5176 12256 5188
rect 12308 5176 12314 5228
rect 12526 5176 12532 5228
rect 12584 5216 12590 5228
rect 12621 5219 12679 5225
rect 12621 5216 12633 5219
rect 12584 5188 12633 5216
rect 12584 5176 12590 5188
rect 12621 5185 12633 5188
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 14826 5176 14832 5228
rect 14884 5176 14890 5228
rect 15028 5225 15056 5256
rect 15470 5244 15476 5256
rect 15528 5244 15534 5296
rect 16132 5284 16160 5312
rect 16850 5284 16856 5296
rect 15856 5256 16856 5284
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5185 15071 5219
rect 15013 5179 15071 5185
rect 15194 5176 15200 5228
rect 15252 5176 15258 5228
rect 15856 5225 15884 5256
rect 16850 5244 16856 5256
rect 16908 5244 16914 5296
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16022 5216 16028 5228
rect 15979 5188 16028 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16022 5176 16028 5188
rect 16080 5176 16086 5228
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 17126 5216 17132 5228
rect 16163 5188 17132 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 17126 5176 17132 5188
rect 17184 5176 17190 5228
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12544 5120 12909 5148
rect 12544 5089 12572 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 14921 5151 14979 5157
rect 14921 5117 14933 5151
rect 14967 5148 14979 5151
rect 16206 5148 16212 5160
rect 14967 5120 16212 5148
rect 14967 5117 14979 5120
rect 14921 5111 14979 5117
rect 16206 5108 16212 5120
rect 16264 5108 16270 5160
rect 12529 5083 12587 5089
rect 10275 5052 10548 5080
rect 12360 5052 12480 5080
rect 10275 5049 10287 5052
rect 10229 5043 10287 5049
rect 4617 5015 4675 5021
rect 4617 4981 4629 5015
rect 4663 5012 4675 5015
rect 4706 5012 4712 5024
rect 4663 4984 4712 5012
rect 4663 4981 4675 4984
rect 4617 4975 4675 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5077 5015 5135 5021
rect 5077 4981 5089 5015
rect 5123 5012 5135 5015
rect 5258 5012 5264 5024
rect 5123 4984 5264 5012
rect 5123 4981 5135 4984
rect 5077 4975 5135 4981
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 12360 5021 12388 5052
rect 12345 5015 12403 5021
rect 12345 4981 12357 5015
rect 12391 4981 12403 5015
rect 12452 5012 12480 5052
rect 12529 5049 12541 5083
rect 12575 5049 12587 5083
rect 12529 5043 12587 5049
rect 15749 5083 15807 5089
rect 15749 5049 15761 5083
rect 15795 5080 15807 5083
rect 16298 5080 16304 5092
rect 15795 5052 16304 5080
rect 15795 5049 15807 5052
rect 15749 5043 15807 5049
rect 16298 5040 16304 5052
rect 16356 5040 16362 5092
rect 14458 5012 14464 5024
rect 12452 4984 14464 5012
rect 12345 4975 12403 4981
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 15562 4972 15568 5024
rect 15620 4972 15626 5024
rect 1104 4922 18860 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 18860 4922
rect 1104 4848 18860 4870
rect 5534 4768 5540 4820
rect 5592 4808 5598 4820
rect 5902 4808 5908 4820
rect 5592 4780 5908 4808
rect 5592 4768 5598 4780
rect 5902 4768 5908 4780
rect 5960 4808 5966 4820
rect 6638 4808 6644 4820
rect 5960 4780 6644 4808
rect 5960 4768 5966 4780
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 9030 4768 9036 4820
rect 9088 4768 9094 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 9493 4811 9551 4817
rect 9493 4808 9505 4811
rect 9364 4780 9505 4808
rect 9364 4768 9370 4780
rect 9493 4777 9505 4780
rect 9539 4777 9551 4811
rect 9493 4771 9551 4777
rect 13630 4768 13636 4820
rect 13688 4768 13694 4820
rect 9398 4740 9404 4752
rect 9048 4712 9404 4740
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 4522 4672 4528 4684
rect 4203 4644 4528 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 4522 4632 4528 4644
rect 4580 4632 4586 4684
rect 9048 4672 9076 4712
rect 9398 4700 9404 4712
rect 9456 4700 9462 4752
rect 8956 4644 9076 4672
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 5810 4564 5816 4616
rect 5868 4604 5874 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 5868 4576 6745 4604
rect 5868 4564 5874 4576
rect 6733 4573 6745 4576
rect 6779 4604 6791 4607
rect 6822 4604 6828 4616
rect 6779 4576 6828 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 6822 4564 6828 4576
rect 6880 4604 6886 4616
rect 8754 4604 8760 4616
rect 6880 4576 8760 4604
rect 6880 4564 6886 4576
rect 8754 4564 8760 4576
rect 8812 4564 8818 4616
rect 8956 4613 8984 4644
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9180 4644 9352 4672
rect 9180 4632 9186 4644
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 9030 4564 9036 4616
rect 9088 4604 9094 4616
rect 9324 4613 9352 4644
rect 9217 4607 9275 4613
rect 9217 4604 9229 4607
rect 9088 4576 9229 4604
rect 9088 4564 9094 4576
rect 9217 4573 9229 4576
rect 9263 4573 9275 4607
rect 9217 4567 9275 4573
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 12342 4564 12348 4616
rect 12400 4604 12406 4616
rect 12437 4607 12495 4613
rect 12437 4604 12449 4607
rect 12400 4576 12449 4604
rect 12400 4564 12406 4576
rect 12437 4573 12449 4576
rect 12483 4573 12495 4607
rect 12437 4567 12495 4573
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 12676 4576 13553 4604
rect 12676 4564 12682 4576
rect 13541 4573 13553 4576
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 4430 4496 4436 4548
rect 4488 4496 4494 4548
rect 6638 4496 6644 4548
rect 6696 4496 6702 4548
rect 6917 4539 6975 4545
rect 6917 4505 6929 4539
rect 6963 4536 6975 4539
rect 9048 4536 9076 4564
rect 6963 4508 9076 4536
rect 6963 4505 6975 4508
rect 6917 4499 6975 4505
rect 6362 4428 6368 4480
rect 6420 4428 6426 4480
rect 6454 4428 6460 4480
rect 6512 4468 6518 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 6512 4440 6561 4468
rect 6512 4428 6518 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6549 4431 6607 4437
rect 12342 4428 12348 4480
rect 12400 4428 12406 4480
rect 1104 4378 18860 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 18860 4378
rect 1104 4304 18860 4326
rect 4430 4224 4436 4276
rect 4488 4264 4494 4276
rect 4525 4267 4583 4273
rect 4525 4264 4537 4267
rect 4488 4236 4537 4264
rect 4488 4224 4494 4236
rect 4525 4233 4537 4236
rect 4571 4233 4583 4267
rect 4525 4227 4583 4233
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 8297 4267 8355 4273
rect 4672 4236 6592 4264
rect 4672 4224 4678 4236
rect 4706 4156 4712 4208
rect 4764 4156 4770 4208
rect 5537 4199 5595 4205
rect 5537 4165 5549 4199
rect 5583 4196 5595 4199
rect 5810 4196 5816 4208
rect 5583 4168 5816 4196
rect 5583 4165 5595 4168
rect 5537 4159 5595 4165
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 6043 4165 6101 4171
rect 5077 4131 5135 4137
rect 5077 4097 5089 4131
rect 5123 4128 5135 4131
rect 5258 4128 5264 4140
rect 5123 4100 5264 4128
rect 5123 4097 5135 4100
rect 5077 4091 5135 4097
rect 5258 4088 5264 4100
rect 5316 4128 5322 4140
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 5316 4100 5365 4128
rect 5316 4088 5322 4100
rect 5353 4097 5365 4100
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 6043 4131 6055 4165
rect 6089 4131 6101 4165
rect 6564 4140 6592 4236
rect 8297 4233 8309 4267
rect 8343 4264 8355 4267
rect 8754 4264 8760 4276
rect 8343 4236 8760 4264
rect 8343 4233 8355 4236
rect 8297 4227 8355 4233
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 9398 4224 9404 4276
rect 9456 4264 9462 4276
rect 11701 4267 11759 4273
rect 11701 4264 11713 4267
rect 9456 4236 11713 4264
rect 9456 4224 9462 4236
rect 11701 4233 11713 4236
rect 11747 4233 11759 4267
rect 11701 4227 11759 4233
rect 12069 4267 12127 4273
rect 12069 4233 12081 4267
rect 12115 4264 12127 4267
rect 12250 4264 12256 4276
rect 12115 4236 12256 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 8050 4168 8524 4196
rect 6043 4128 6101 4131
rect 6454 4128 6460 4140
rect 5500 4100 6460 4128
rect 5500 4088 5506 4100
rect 6454 4088 6460 4100
rect 6512 4088 6518 4140
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 8496 4137 8524 4168
rect 10502 4156 10508 4208
rect 10560 4156 10566 4208
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 11793 4199 11851 4205
rect 11793 4196 11805 4199
rect 11112 4168 11805 4196
rect 11112 4156 11118 4168
rect 11793 4165 11805 4168
rect 11839 4165 11851 4199
rect 11793 4159 11851 4165
rect 13814 4156 13820 4208
rect 13872 4156 13878 4208
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4097 8539 4131
rect 8481 4091 8539 4097
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 9214 4128 9220 4140
rect 8619 4100 9220 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 9950 4128 9956 4140
rect 9732 4100 9956 4128
rect 9732 4088 9738 4100
rect 9950 4088 9956 4100
rect 10008 4128 10014 4140
rect 10686 4128 10692 4140
rect 10008 4100 10692 4128
rect 10008 4088 10014 4100
rect 10686 4088 10692 4100
rect 10744 4128 10750 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 10744 4100 11529 4128
rect 10744 4088 10750 4100
rect 11517 4097 11529 4100
rect 11563 4128 11575 4131
rect 11698 4128 11704 4140
rect 11563 4100 11704 4128
rect 11563 4097 11575 4100
rect 11517 4091 11575 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 12158 4128 12164 4140
rect 11992 4100 12164 4128
rect 6822 4020 6828 4072
rect 6880 4020 6886 4072
rect 8202 4020 8208 4072
rect 8260 4060 8266 4072
rect 11992 4060 12020 4100
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12342 4088 12348 4140
rect 12400 4088 12406 4140
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 8260 4032 12020 4060
rect 8260 4020 8266 4032
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12452 4060 12480 4091
rect 12124 4032 12480 4060
rect 12124 4020 12130 4032
rect 10134 3952 10140 4004
rect 10192 3952 10198 4004
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 10689 3995 10747 4001
rect 10689 3992 10701 3995
rect 10468 3964 10701 3992
rect 10468 3952 10474 3964
rect 10689 3961 10701 3964
rect 10735 3961 10747 3995
rect 12544 3992 12572 4091
rect 12618 4088 12624 4140
rect 12676 4128 12682 4140
rect 12897 4131 12955 4137
rect 12897 4128 12909 4131
rect 12676 4100 12909 4128
rect 12676 4088 12682 4100
rect 12897 4097 12909 4100
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12805 4063 12863 4069
rect 12805 4029 12817 4063
rect 12851 4060 12863 4063
rect 13173 4063 13231 4069
rect 13173 4060 13185 4063
rect 12851 4032 13185 4060
rect 12851 4029 12863 4032
rect 12805 4023 12863 4029
rect 13173 4029 13185 4032
rect 13219 4029 13231 4063
rect 13173 4023 13231 4029
rect 12618 3992 12624 4004
rect 12544 3964 12624 3992
rect 10689 3955 10747 3961
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 4798 3924 4804 3936
rect 4755 3896 4804 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5718 3884 5724 3936
rect 5776 3884 5782 3936
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5960 3896 6009 3924
rect 5960 3884 5966 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 5997 3887 6055 3893
rect 6178 3884 6184 3936
rect 6236 3884 6242 3936
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10594 3924 10600 3936
rect 10551 3896 10600 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10594 3884 10600 3896
rect 10652 3884 10658 3936
rect 12636 3924 12664 3952
rect 14550 3924 14556 3936
rect 12636 3896 14556 3924
rect 14550 3884 14556 3896
rect 14608 3924 14614 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 14608 3896 14657 3924
rect 14608 3884 14614 3896
rect 14645 3893 14657 3896
rect 14691 3893 14703 3927
rect 14645 3887 14703 3893
rect 1104 3834 18860 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 18860 3834
rect 1104 3760 18860 3782
rect 5169 3723 5227 3729
rect 5169 3689 5181 3723
rect 5215 3720 5227 3723
rect 5534 3720 5540 3732
rect 5215 3692 5540 3720
rect 5215 3689 5227 3692
rect 5169 3683 5227 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 6104 3692 6561 3720
rect 4798 3612 4804 3664
rect 4856 3652 4862 3664
rect 6104 3652 6132 3692
rect 6549 3689 6561 3692
rect 6595 3689 6607 3723
rect 6549 3683 6607 3689
rect 6733 3723 6791 3729
rect 6733 3689 6745 3723
rect 6779 3720 6791 3723
rect 6822 3720 6828 3732
rect 6779 3692 6828 3720
rect 6779 3689 6791 3692
rect 6733 3683 6791 3689
rect 4856 3624 6132 3652
rect 4856 3612 4862 3624
rect 6178 3612 6184 3664
rect 6236 3612 6242 3664
rect 6564 3652 6592 3683
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 9493 3723 9551 3729
rect 9493 3720 9505 3723
rect 8619 3692 9505 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 9493 3689 9505 3692
rect 9539 3689 9551 3723
rect 9861 3723 9919 3729
rect 9861 3720 9873 3723
rect 9493 3683 9551 3689
rect 9646 3692 9873 3720
rect 7006 3652 7012 3664
rect 6564 3624 7012 3652
rect 7006 3612 7012 3624
rect 7064 3652 7070 3664
rect 8202 3652 8208 3664
rect 7064 3624 8208 3652
rect 7064 3612 7070 3624
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 9398 3612 9404 3664
rect 9456 3652 9462 3664
rect 9646 3652 9674 3692
rect 9861 3689 9873 3692
rect 9907 3689 9919 3723
rect 9861 3683 9919 3689
rect 10045 3723 10103 3729
rect 10045 3689 10057 3723
rect 10091 3720 10103 3723
rect 10134 3720 10140 3732
rect 10091 3692 10140 3720
rect 10091 3689 10103 3692
rect 10045 3683 10103 3689
rect 10134 3680 10140 3692
rect 10192 3720 10198 3732
rect 10192 3692 11468 3720
rect 10192 3680 10198 3692
rect 9456 3624 9674 3652
rect 11440 3652 11468 3692
rect 11882 3680 11888 3732
rect 11940 3720 11946 3732
rect 12253 3723 12311 3729
rect 12253 3720 12265 3723
rect 11940 3692 12265 3720
rect 11940 3680 11946 3692
rect 12253 3689 12265 3692
rect 12299 3689 12311 3723
rect 12253 3683 12311 3689
rect 12342 3680 12348 3732
rect 12400 3720 12406 3732
rect 12400 3692 13768 3720
rect 12400 3680 12406 3692
rect 11440 3624 12434 3652
rect 9456 3612 9462 3624
rect 5261 3519 5319 3525
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 6196 3516 6224 3612
rect 6362 3544 6368 3596
rect 6420 3584 6426 3596
rect 6420 3556 9628 3584
rect 6420 3544 6426 3556
rect 6825 3519 6883 3525
rect 6825 3516 6837 3519
rect 5307 3488 5672 3516
rect 6196 3488 6837 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 5644 3380 5672 3488
rect 6825 3485 6837 3488
rect 6871 3485 6883 3519
rect 6825 3479 6883 3485
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3516 7067 3519
rect 8846 3516 8852 3528
rect 7055 3488 8852 3516
rect 7055 3485 7067 3488
rect 7009 3479 7067 3485
rect 8846 3476 8852 3488
rect 8904 3476 8910 3528
rect 9324 3525 9352 3556
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 9398 3476 9404 3528
rect 9456 3476 9462 3528
rect 9600 3525 9628 3556
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 11698 3544 11704 3596
rect 11756 3584 11762 3596
rect 11885 3587 11943 3593
rect 11885 3584 11897 3587
rect 11756 3556 11897 3584
rect 11756 3544 11762 3556
rect 11885 3553 11897 3556
rect 11931 3553 11943 3587
rect 12406 3584 12434 3624
rect 12406 3556 13216 3584
rect 11885 3547 11943 3553
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3516 9643 3519
rect 9631 3488 9812 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 5718 3408 5724 3460
rect 5776 3448 5782 3460
rect 6549 3451 6607 3457
rect 6549 3448 6561 3451
rect 5776 3420 6561 3448
rect 5776 3408 5782 3420
rect 6549 3417 6561 3420
rect 6595 3417 6607 3451
rect 6914 3448 6920 3460
rect 6549 3411 6607 3417
rect 6656 3420 6920 3448
rect 6656 3380 6684 3420
rect 6914 3408 6920 3420
rect 6972 3448 6978 3460
rect 8110 3448 8116 3460
rect 6972 3420 8116 3448
rect 6972 3408 6978 3420
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8202 3408 8208 3460
rect 8260 3448 8266 3460
rect 8389 3451 8447 3457
rect 8389 3448 8401 3451
rect 8260 3420 8401 3448
rect 8260 3408 8266 3420
rect 8389 3417 8401 3420
rect 8435 3417 8447 3451
rect 8389 3411 8447 3417
rect 8605 3451 8663 3457
rect 8605 3417 8617 3451
rect 8651 3448 8663 3451
rect 8941 3451 8999 3457
rect 8941 3448 8953 3451
rect 8651 3420 8953 3448
rect 8651 3417 8663 3420
rect 8605 3411 8663 3417
rect 8941 3417 8953 3420
rect 8987 3417 8999 3451
rect 8941 3411 8999 3417
rect 9125 3451 9183 3457
rect 9125 3417 9137 3451
rect 9171 3448 9183 3451
rect 9416 3448 9444 3476
rect 9171 3420 9444 3448
rect 9171 3417 9183 3420
rect 9125 3411 9183 3417
rect 9674 3408 9680 3460
rect 9732 3408 9738 3460
rect 9784 3448 9812 3488
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 11514 3476 11520 3528
rect 11572 3476 11578 3528
rect 12437 3519 12495 3525
rect 12437 3485 12449 3519
rect 12483 3485 12495 3519
rect 12437 3479 12495 3485
rect 9877 3451 9935 3457
rect 9877 3448 9889 3451
rect 9784 3420 9889 3448
rect 9877 3417 9889 3420
rect 9923 3448 9935 3451
rect 12452 3448 12480 3479
rect 12618 3476 12624 3528
rect 12676 3476 12682 3528
rect 12912 3525 12940 3556
rect 13188 3525 13216 3556
rect 12897 3519 12955 3525
rect 12897 3485 12909 3519
rect 12943 3485 12955 3519
rect 12897 3479 12955 3485
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 13096 3448 13124 3479
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 13740 3525 13768 3692
rect 13814 3680 13820 3732
rect 13872 3680 13878 3732
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13688 3488 13737 3516
rect 13688 3476 13694 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 13357 3451 13415 3457
rect 13357 3448 13369 3451
rect 9923 3420 10824 3448
rect 12452 3420 13369 3448
rect 9923 3417 9935 3420
rect 9877 3411 9935 3417
rect 5644 3352 6684 3380
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 8757 3383 8815 3389
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 8846 3380 8852 3392
rect 8803 3352 8852 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 10796 3380 10824 3420
rect 13357 3417 13369 3420
rect 13403 3448 13415 3451
rect 14826 3448 14832 3460
rect 13403 3420 14832 3448
rect 13403 3417 13415 3420
rect 13357 3411 13415 3417
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 11054 3380 11060 3392
rect 10796 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 12066 3340 12072 3392
rect 12124 3380 12130 3392
rect 12713 3383 12771 3389
rect 12713 3380 12725 3383
rect 12124 3352 12725 3380
rect 12124 3340 12130 3352
rect 12713 3349 12725 3352
rect 12759 3349 12771 3383
rect 12713 3343 12771 3349
rect 13538 3340 13544 3392
rect 13596 3340 13602 3392
rect 1104 3290 18860 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 18860 3290
rect 1104 3216 18860 3238
rect 10134 3176 10140 3188
rect 8588 3148 10140 3176
rect 8018 3068 8024 3120
rect 8076 3068 8082 3120
rect 6546 3000 6552 3052
rect 6604 3040 6610 3052
rect 8588 3049 8616 3148
rect 10134 3136 10140 3148
rect 10192 3176 10198 3188
rect 12526 3176 12532 3188
rect 10192 3148 12532 3176
rect 10192 3136 10198 3148
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 14461 3179 14519 3185
rect 14461 3145 14473 3179
rect 14507 3176 14519 3179
rect 14826 3176 14832 3188
rect 14507 3148 14832 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 14826 3136 14832 3148
rect 14884 3136 14890 3188
rect 8846 3068 8852 3120
rect 8904 3068 8910 3120
rect 10410 3108 10416 3120
rect 10074 3080 10416 3108
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 10502 3068 10508 3120
rect 10560 3068 10566 3120
rect 10628 3080 11284 3108
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6604 3012 6745 3040
rect 6604 3000 6610 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3009 8631 3043
rect 8573 3003 8631 3009
rect 7009 2975 7067 2981
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7098 2972 7104 2984
rect 7055 2944 7104 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 8481 2975 8539 2981
rect 8481 2941 8493 2975
rect 8527 2972 8539 2975
rect 8938 2972 8944 2984
rect 8527 2944 8944 2972
rect 8527 2941 8539 2944
rect 8481 2935 8539 2941
rect 8938 2932 8944 2944
rect 8996 2932 9002 2984
rect 9214 2932 9220 2984
rect 9272 2972 9278 2984
rect 10628 2972 10656 3080
rect 10686 3000 10692 3052
rect 10744 3000 10750 3052
rect 10873 3043 10931 3049
rect 10873 3040 10885 3043
rect 10796 3012 10885 3040
rect 9272 2944 10656 2972
rect 9272 2932 9278 2944
rect 10321 2907 10379 2913
rect 10321 2873 10333 2907
rect 10367 2904 10379 2907
rect 10796 2904 10824 3012
rect 10873 3009 10885 3012
rect 10919 3009 10931 3043
rect 10873 3003 10931 3009
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3040 11023 3043
rect 11054 3040 11060 3052
rect 11011 3012 11060 3040
rect 11011 3009 11023 3012
rect 10965 3003 11023 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11256 3049 11284 3080
rect 11514 3068 11520 3120
rect 11572 3108 11578 3120
rect 11609 3111 11667 3117
rect 11609 3108 11621 3111
rect 11572 3080 11621 3108
rect 11572 3068 11578 3080
rect 11609 3077 11621 3080
rect 11655 3077 11667 3111
rect 12342 3108 12348 3120
rect 11609 3071 11667 3077
rect 11716 3080 12348 3108
rect 11716 3049 11744 3080
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3077 12495 3111
rect 12437 3071 12495 3077
rect 11241 3043 11299 3049
rect 11241 3009 11253 3043
rect 11287 3040 11299 3043
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11287 3012 11713 3040
rect 11287 3009 11299 3012
rect 11241 3003 11299 3009
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11701 3003 11759 3009
rect 12066 3000 12072 3052
rect 12124 3000 12130 3052
rect 12452 2904 12480 3071
rect 12544 3040 12572 3136
rect 13998 3068 14004 3120
rect 14056 3068 14062 3120
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12544 3012 12725 3040
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12713 3003 12771 3009
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12636 2944 13001 2972
rect 12636 2913 12664 2944
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 12989 2935 13047 2941
rect 10367 2876 10824 2904
rect 10980 2876 12480 2904
rect 12621 2907 12679 2913
rect 10367 2873 10379 2876
rect 10321 2867 10379 2873
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 9214 2836 9220 2848
rect 8168 2808 9220 2836
rect 8168 2796 8174 2808
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 10336 2836 10364 2867
rect 9456 2808 10364 2836
rect 9456 2796 9462 2808
rect 10594 2796 10600 2848
rect 10652 2836 10658 2848
rect 10980 2836 11008 2876
rect 12621 2873 12633 2907
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 10652 2808 11008 2836
rect 12437 2839 12495 2845
rect 10652 2796 10658 2808
rect 12437 2805 12449 2839
rect 12483 2836 12495 2839
rect 13538 2836 13544 2848
rect 12483 2808 13544 2836
rect 12483 2805 12495 2808
rect 12437 2799 12495 2805
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 1104 2746 18860 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 18860 2746
rect 1104 2672 18860 2694
rect 7006 2592 7012 2644
rect 7064 2592 7070 2644
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7193 2635 7251 2641
rect 7193 2632 7205 2635
rect 7156 2604 7205 2632
rect 7156 2592 7162 2604
rect 7193 2601 7205 2604
rect 7239 2601 7251 2635
rect 7193 2595 7251 2601
rect 8018 2592 8024 2644
rect 8076 2592 8082 2644
rect 8662 2592 8668 2644
rect 8720 2592 8726 2644
rect 13725 2635 13783 2641
rect 13725 2601 13737 2635
rect 13771 2632 13783 2635
rect 13998 2632 14004 2644
rect 13771 2604 14004 2632
rect 13771 2601 13783 2604
rect 13725 2595 13783 2601
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 6362 2524 6368 2576
rect 6420 2564 6426 2576
rect 6641 2567 6699 2573
rect 6641 2564 6653 2567
rect 6420 2536 6653 2564
rect 6420 2524 6426 2536
rect 6641 2533 6653 2536
rect 6687 2533 6699 2567
rect 6641 2527 6699 2533
rect 8478 2524 8484 2576
rect 8536 2564 8542 2576
rect 9401 2567 9459 2573
rect 9401 2564 9413 2567
rect 8536 2536 9413 2564
rect 8536 2524 8542 2536
rect 9401 2533 9413 2536
rect 9447 2533 9459 2567
rect 9401 2527 9459 2533
rect 9766 2524 9772 2576
rect 9824 2564 9830 2576
rect 9824 2536 10088 2564
rect 9824 2524 9830 2536
rect 10060 2505 10088 2536
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2465 10103 2499
rect 10045 2459 10103 2465
rect 8110 2388 8116 2440
rect 8168 2388 8174 2440
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 7009 2363 7067 2369
rect 7009 2329 7021 2363
rect 7055 2360 7067 2363
rect 7190 2360 7196 2372
rect 7055 2332 7196 2360
rect 7055 2329 7067 2332
rect 7009 2323 7067 2329
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 7742 2320 7748 2372
rect 7800 2360 7806 2372
rect 8220 2360 8248 2391
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8444 2400 8493 2428
rect 8444 2388 8450 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 13630 2388 13636 2440
rect 13688 2388 13694 2440
rect 7800 2332 8248 2360
rect 7800 2320 7806 2332
rect 9030 2320 9036 2372
rect 9088 2360 9094 2372
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 9088 2332 9229 2360
rect 9088 2320 9094 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 8389 2295 8447 2301
rect 8389 2261 8401 2295
rect 8435 2292 8447 2295
rect 8754 2292 8760 2304
rect 8435 2264 8760 2292
rect 8435 2261 8447 2264
rect 8389 2255 8447 2261
rect 8754 2252 8760 2264
rect 8812 2252 8818 2304
rect 1104 2202 18860 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 18860 2202
rect 1104 2128 18860 2150
<< via1 >>
rect 14832 20680 14884 20732
rect 16856 20680 16908 20732
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 14188 19456 14240 19508
rect 15936 19456 15988 19508
rect 7012 19388 7064 19440
rect 5632 19184 5684 19236
rect 6092 19363 6144 19372
rect 6092 19329 6101 19363
rect 6101 19329 6135 19363
rect 6135 19329 6144 19363
rect 6092 19320 6144 19329
rect 6184 19363 6236 19372
rect 6184 19329 6193 19363
rect 6193 19329 6227 19363
rect 6227 19329 6236 19363
rect 6184 19320 6236 19329
rect 6460 19320 6512 19372
rect 11336 19320 11388 19372
rect 13268 19363 13320 19372
rect 13268 19329 13277 19363
rect 13277 19329 13311 19363
rect 13311 19329 13320 19363
rect 13268 19320 13320 19329
rect 14188 19363 14240 19372
rect 14188 19329 14197 19363
rect 14197 19329 14231 19363
rect 14231 19329 14240 19363
rect 14188 19320 14240 19329
rect 15936 19363 15988 19372
rect 15936 19329 15945 19363
rect 15945 19329 15979 19363
rect 15979 19329 15988 19363
rect 15936 19320 15988 19329
rect 5816 19252 5868 19304
rect 6644 19295 6696 19304
rect 6644 19261 6653 19295
rect 6653 19261 6687 19295
rect 6687 19261 6696 19295
rect 6644 19252 6696 19261
rect 12900 19252 12952 19304
rect 9312 19184 9364 19236
rect 14280 19184 14332 19236
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 15476 19295 15528 19304
rect 15476 19261 15485 19295
rect 15485 19261 15519 19295
rect 15519 19261 15528 19295
rect 15476 19252 15528 19261
rect 16120 19227 16172 19236
rect 16120 19193 16129 19227
rect 16129 19193 16163 19227
rect 16163 19193 16172 19227
rect 16120 19184 16172 19193
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 11244 19116 11296 19168
rect 14372 19159 14424 19168
rect 14372 19125 14381 19159
rect 14381 19125 14415 19159
rect 14415 19125 14424 19159
rect 14372 19116 14424 19125
rect 14832 19116 14884 19168
rect 16488 19184 16540 19236
rect 16304 19159 16356 19168
rect 16304 19125 16313 19159
rect 16313 19125 16347 19159
rect 16347 19125 16356 19159
rect 16304 19116 16356 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 4620 18751 4672 18760
rect 4620 18717 4629 18751
rect 4629 18717 4663 18751
rect 4663 18717 4672 18751
rect 4620 18708 4672 18717
rect 5816 18912 5868 18964
rect 9864 18912 9916 18964
rect 11336 18912 11388 18964
rect 5724 18776 5776 18828
rect 10784 18776 10836 18828
rect 15384 18912 15436 18964
rect 16120 18887 16172 18896
rect 16120 18853 16129 18887
rect 16129 18853 16163 18887
rect 16163 18853 16172 18887
rect 16120 18844 16172 18853
rect 4344 18640 4396 18692
rect 6460 18708 6512 18760
rect 14188 18751 14240 18760
rect 14188 18717 14197 18751
rect 14197 18717 14231 18751
rect 14231 18717 14240 18751
rect 14188 18708 14240 18717
rect 14280 18708 14332 18760
rect 14832 18751 14884 18760
rect 14832 18717 14841 18751
rect 14841 18717 14875 18751
rect 14875 18717 14884 18751
rect 14832 18708 14884 18717
rect 4620 18572 4672 18624
rect 5264 18640 5316 18692
rect 10232 18683 10284 18692
rect 10232 18649 10241 18683
rect 10241 18649 10275 18683
rect 10275 18649 10284 18683
rect 10232 18640 10284 18649
rect 11244 18640 11296 18692
rect 12072 18683 12124 18692
rect 12072 18649 12081 18683
rect 12081 18649 12115 18683
rect 12115 18649 12124 18683
rect 12072 18640 12124 18649
rect 15936 18776 15988 18828
rect 15292 18683 15344 18692
rect 15292 18649 15301 18683
rect 15301 18649 15335 18683
rect 15335 18649 15344 18683
rect 15292 18640 15344 18649
rect 6736 18572 6788 18624
rect 11704 18615 11756 18624
rect 11704 18581 11713 18615
rect 11713 18581 11747 18615
rect 11747 18581 11756 18615
rect 11704 18572 11756 18581
rect 13084 18572 13136 18624
rect 13544 18615 13596 18624
rect 13544 18581 13553 18615
rect 13553 18581 13587 18615
rect 13587 18581 13596 18615
rect 13544 18572 13596 18581
rect 13728 18572 13780 18624
rect 16304 18708 16356 18760
rect 16488 18708 16540 18760
rect 15752 18615 15804 18624
rect 15752 18581 15761 18615
rect 15761 18581 15795 18615
rect 15795 18581 15804 18615
rect 15752 18572 15804 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 5632 18368 5684 18420
rect 6460 18411 6512 18420
rect 6460 18377 6469 18411
rect 6469 18377 6503 18411
rect 6503 18377 6512 18411
rect 6460 18368 6512 18377
rect 10232 18368 10284 18420
rect 12072 18411 12124 18420
rect 12072 18377 12081 18411
rect 12081 18377 12115 18411
rect 12115 18377 12124 18411
rect 12072 18368 12124 18377
rect 4620 18343 4672 18352
rect 4620 18309 4629 18343
rect 4629 18309 4663 18343
rect 4663 18309 4672 18343
rect 4620 18300 4672 18309
rect 6092 18300 6144 18352
rect 4344 18275 4396 18284
rect 4344 18241 4353 18275
rect 4353 18241 4387 18275
rect 4387 18241 4396 18275
rect 4344 18232 4396 18241
rect 6184 18232 6236 18284
rect 7748 18232 7800 18284
rect 9864 18232 9916 18284
rect 11520 18300 11572 18352
rect 11888 18343 11940 18352
rect 11888 18309 11897 18343
rect 11897 18309 11931 18343
rect 11931 18309 11940 18343
rect 11888 18300 11940 18309
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 11152 18232 11204 18284
rect 13084 18368 13136 18420
rect 13452 18368 13504 18420
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 14372 18368 14424 18420
rect 15016 18368 15068 18420
rect 12900 18300 12952 18352
rect 15476 18300 15528 18352
rect 5356 18164 5408 18216
rect 11704 18164 11756 18216
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 13820 18232 13872 18284
rect 14832 18232 14884 18284
rect 15292 18232 15344 18284
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 13452 18096 13504 18148
rect 15936 18096 15988 18148
rect 4712 18028 4764 18080
rect 5356 18028 5408 18080
rect 9496 18071 9548 18080
rect 9496 18037 9505 18071
rect 9505 18037 9539 18071
rect 9539 18037 9548 18071
rect 9496 18028 9548 18037
rect 11244 18028 11296 18080
rect 12256 18071 12308 18080
rect 12256 18037 12265 18071
rect 12265 18037 12299 18071
rect 12299 18037 12308 18071
rect 12256 18028 12308 18037
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 13544 18028 13596 18080
rect 15568 18028 15620 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2596 17867 2648 17876
rect 2596 17833 2605 17867
rect 2605 17833 2639 17867
rect 2639 17833 2648 17867
rect 2596 17824 2648 17833
rect 5264 17824 5316 17876
rect 4068 17756 4120 17808
rect 6184 17824 6236 17876
rect 10508 17824 10560 17876
rect 11888 17824 11940 17876
rect 14924 17799 14976 17808
rect 14924 17765 14933 17799
rect 14933 17765 14967 17799
rect 14967 17765 14976 17799
rect 14924 17756 14976 17765
rect 15844 17756 15896 17808
rect 2872 17688 2924 17740
rect 3976 17688 4028 17740
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 5356 17688 5408 17740
rect 10048 17688 10100 17740
rect 10784 17731 10836 17740
rect 10784 17697 10793 17731
rect 10793 17697 10827 17731
rect 10827 17697 10836 17731
rect 10784 17688 10836 17697
rect 6276 17663 6328 17672
rect 6276 17629 6285 17663
rect 6285 17629 6319 17663
rect 6319 17629 6328 17663
rect 6276 17620 6328 17629
rect 2412 17527 2464 17536
rect 2412 17493 2421 17527
rect 2421 17493 2455 17527
rect 2455 17493 2464 17527
rect 2412 17484 2464 17493
rect 2504 17484 2556 17536
rect 9496 17552 9548 17604
rect 5724 17484 5776 17536
rect 6460 17484 6512 17536
rect 7104 17484 7156 17536
rect 10324 17484 10376 17536
rect 10600 17552 10652 17604
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 12256 17620 12308 17672
rect 14188 17620 14240 17672
rect 14832 17620 14884 17672
rect 15752 17688 15804 17740
rect 11152 17552 11204 17604
rect 15016 17552 15068 17604
rect 15476 17620 15528 17672
rect 15568 17663 15620 17672
rect 15568 17629 15577 17663
rect 15577 17629 15611 17663
rect 15611 17629 15620 17663
rect 15568 17620 15620 17629
rect 14280 17484 14332 17536
rect 15292 17484 15344 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2412 17280 2464 17332
rect 3148 17280 3200 17332
rect 4068 17323 4120 17332
rect 4068 17289 4077 17323
rect 4077 17289 4111 17323
rect 4111 17289 4120 17323
rect 4068 17280 4120 17289
rect 5356 17280 5408 17332
rect 6184 17323 6236 17332
rect 6184 17289 6193 17323
rect 6193 17289 6227 17323
rect 6227 17289 6236 17323
rect 6184 17280 6236 17289
rect 7748 17280 7800 17332
rect 1768 17212 1820 17264
rect 2504 17212 2556 17264
rect 2320 17144 2372 17196
rect 3056 17187 3108 17196
rect 3056 17153 3065 17187
rect 3065 17153 3099 17187
rect 3099 17153 3108 17187
rect 3056 17144 3108 17153
rect 3240 17144 3292 17196
rect 3976 17212 4028 17264
rect 7012 17212 7064 17264
rect 7104 17255 7156 17264
rect 7104 17221 7113 17255
rect 7113 17221 7147 17255
rect 7147 17221 7156 17255
rect 7104 17212 7156 17221
rect 4804 17144 4856 17196
rect 5724 17187 5776 17196
rect 5724 17153 5733 17187
rect 5733 17153 5767 17187
rect 5767 17153 5776 17187
rect 5724 17144 5776 17153
rect 6092 17144 6144 17196
rect 6736 17144 6788 17196
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 15108 17280 15160 17332
rect 10324 17255 10376 17264
rect 10324 17221 10333 17255
rect 10333 17221 10367 17255
rect 10367 17221 10376 17255
rect 10324 17212 10376 17221
rect 9312 17144 9364 17196
rect 9956 17144 10008 17196
rect 4620 17076 4672 17128
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 12808 17076 12860 17128
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 12440 17008 12492 17060
rect 1952 16940 2004 16992
rect 2412 16940 2464 16992
rect 3332 16983 3384 16992
rect 3332 16949 3341 16983
rect 3341 16949 3375 16983
rect 3375 16949 3384 16983
rect 3332 16940 3384 16949
rect 4712 16940 4764 16992
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 12716 16983 12768 16992
rect 12716 16949 12725 16983
rect 12725 16949 12759 16983
rect 12759 16949 12768 16983
rect 12716 16940 12768 16949
rect 13084 16940 13136 16992
rect 13728 16940 13780 16992
rect 14648 17187 14700 17196
rect 14648 17153 14657 17187
rect 14657 17153 14691 17187
rect 14691 17153 14700 17187
rect 14648 17144 14700 17153
rect 14740 17187 14792 17196
rect 14740 17153 14749 17187
rect 14749 17153 14783 17187
rect 14783 17153 14792 17187
rect 14740 17144 14792 17153
rect 14832 17187 14884 17196
rect 14832 17153 14841 17187
rect 14841 17153 14875 17187
rect 14875 17153 14884 17187
rect 14832 17144 14884 17153
rect 15016 17187 15068 17196
rect 15016 17153 15025 17187
rect 15025 17153 15059 17187
rect 15059 17153 15068 17187
rect 15016 17144 15068 17153
rect 15936 17144 15988 17196
rect 15476 17076 15528 17128
rect 15568 17008 15620 17060
rect 15844 17008 15896 17060
rect 15016 16940 15068 16992
rect 15384 16983 15436 16992
rect 15384 16949 15393 16983
rect 15393 16949 15427 16983
rect 15427 16949 15436 16983
rect 15384 16940 15436 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 2596 16736 2648 16788
rect 3148 16736 3200 16788
rect 1676 16464 1728 16516
rect 1952 16575 2004 16584
rect 1952 16541 1961 16575
rect 1961 16541 1995 16575
rect 1995 16541 2004 16575
rect 1952 16532 2004 16541
rect 2872 16532 2924 16584
rect 2780 16507 2832 16516
rect 2780 16473 2789 16507
rect 2789 16473 2823 16507
rect 2823 16473 2832 16507
rect 2780 16464 2832 16473
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 5540 16736 5592 16788
rect 6276 16736 6328 16788
rect 10416 16779 10468 16788
rect 10416 16745 10425 16779
rect 10425 16745 10459 16779
rect 10459 16745 10468 16779
rect 10416 16736 10468 16745
rect 13728 16779 13780 16788
rect 13728 16745 13737 16779
rect 13737 16745 13771 16779
rect 13771 16745 13780 16779
rect 13728 16736 13780 16745
rect 14372 16736 14424 16788
rect 5356 16668 5408 16720
rect 6644 16600 6696 16652
rect 12808 16600 12860 16652
rect 13360 16600 13412 16652
rect 4620 16532 4672 16541
rect 5356 16532 5408 16584
rect 5724 16532 5776 16584
rect 6000 16532 6052 16584
rect 1860 16439 1912 16448
rect 1860 16405 1869 16439
rect 1869 16405 1903 16439
rect 1903 16405 1912 16439
rect 1860 16396 1912 16405
rect 2596 16396 2648 16448
rect 6276 16532 6328 16584
rect 9128 16464 9180 16516
rect 11980 16532 12032 16584
rect 4620 16439 4672 16448
rect 4620 16405 4629 16439
rect 4629 16405 4663 16439
rect 4663 16405 4672 16439
rect 4620 16396 4672 16405
rect 5356 16396 5408 16448
rect 6000 16439 6052 16448
rect 6000 16405 6009 16439
rect 6009 16405 6043 16439
rect 6043 16405 6052 16439
rect 6000 16396 6052 16405
rect 6092 16439 6144 16448
rect 6092 16405 6101 16439
rect 6101 16405 6135 16439
rect 6135 16405 6144 16439
rect 6092 16396 6144 16405
rect 6276 16439 6328 16448
rect 6276 16405 6285 16439
rect 6285 16405 6319 16439
rect 6319 16405 6328 16439
rect 6276 16396 6328 16405
rect 6644 16396 6696 16448
rect 9956 16396 10008 16448
rect 12440 16507 12492 16516
rect 12440 16473 12449 16507
rect 12449 16473 12483 16507
rect 12483 16473 12492 16507
rect 12440 16464 12492 16473
rect 10876 16396 10928 16448
rect 12992 16439 13044 16448
rect 12992 16405 13001 16439
rect 13001 16405 13035 16439
rect 13035 16405 13044 16439
rect 12992 16396 13044 16405
rect 13176 16439 13228 16448
rect 13176 16405 13185 16439
rect 13185 16405 13219 16439
rect 13219 16405 13228 16439
rect 13176 16396 13228 16405
rect 14556 16600 14608 16652
rect 14280 16575 14332 16584
rect 14280 16541 14289 16575
rect 14289 16541 14323 16575
rect 14323 16541 14332 16575
rect 14280 16532 14332 16541
rect 14924 16575 14976 16584
rect 14924 16541 14933 16575
rect 14933 16541 14967 16575
rect 14967 16541 14976 16575
rect 14924 16532 14976 16541
rect 15476 16575 15528 16584
rect 15476 16541 15485 16575
rect 15485 16541 15519 16575
rect 15519 16541 15528 16575
rect 15476 16532 15528 16541
rect 15568 16532 15620 16584
rect 15844 16532 15896 16584
rect 14372 16396 14424 16448
rect 16212 16396 16264 16448
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 1768 16192 1820 16244
rect 2320 16192 2372 16244
rect 6092 16192 6144 16244
rect 12992 16192 13044 16244
rect 13268 16192 13320 16244
rect 2688 16124 2740 16176
rect 848 16056 900 16108
rect 1860 16056 1912 16108
rect 4804 16124 4856 16176
rect 5356 16124 5408 16176
rect 6460 16124 6512 16176
rect 9036 16124 9088 16176
rect 5724 16056 5776 16108
rect 6276 16056 6328 16108
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 10048 16056 10100 16108
rect 2596 16031 2648 16040
rect 2596 15997 2605 16031
rect 2605 15997 2639 16031
rect 2639 15997 2648 16031
rect 2596 15988 2648 15997
rect 4896 15988 4948 16040
rect 9496 15988 9548 16040
rect 9956 16031 10008 16040
rect 9956 15997 9965 16031
rect 9965 15997 9999 16031
rect 9999 15997 10008 16031
rect 9956 15988 10008 15997
rect 10416 16124 10468 16176
rect 10876 16056 10928 16108
rect 11244 16056 11296 16108
rect 11520 16056 11572 16108
rect 3884 15920 3936 15972
rect 6000 15920 6052 15972
rect 3240 15852 3292 15904
rect 3700 15852 3752 15904
rect 4804 15852 4856 15904
rect 6644 15852 6696 15904
rect 6920 15895 6972 15904
rect 6920 15861 6929 15895
rect 6929 15861 6963 15895
rect 6963 15861 6972 15895
rect 6920 15852 6972 15861
rect 7656 15895 7708 15904
rect 7656 15861 7665 15895
rect 7665 15861 7699 15895
rect 7699 15861 7708 15895
rect 7656 15852 7708 15861
rect 11980 15988 12032 16040
rect 11152 15920 11204 15972
rect 11888 15920 11940 15972
rect 12900 16099 12952 16108
rect 12900 16065 12909 16099
rect 12909 16065 12943 16099
rect 12943 16065 12952 16099
rect 12900 16056 12952 16065
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 14372 16167 14424 16176
rect 14372 16133 14381 16167
rect 14381 16133 14415 16167
rect 14415 16133 14424 16167
rect 14372 16124 14424 16133
rect 14740 16235 14792 16244
rect 14740 16201 14749 16235
rect 14749 16201 14783 16235
rect 14783 16201 14792 16235
rect 14740 16192 14792 16201
rect 16672 16192 16724 16244
rect 13268 16099 13320 16108
rect 13268 16065 13277 16099
rect 13277 16065 13311 16099
rect 13311 16065 13320 16099
rect 13268 16056 13320 16065
rect 13452 16099 13504 16108
rect 13452 16065 13461 16099
rect 13461 16065 13495 16099
rect 13495 16065 13504 16099
rect 13452 16056 13504 16065
rect 14464 16056 14516 16108
rect 15292 16124 15344 16176
rect 15936 16124 15988 16176
rect 14924 16099 14976 16108
rect 14924 16065 14933 16099
rect 14933 16065 14967 16099
rect 14967 16065 14976 16099
rect 14924 16056 14976 16065
rect 15384 16099 15436 16108
rect 15384 16065 15393 16099
rect 15393 16065 15427 16099
rect 15427 16065 15436 16099
rect 15384 16056 15436 16065
rect 16212 16099 16264 16108
rect 16212 16065 16221 16099
rect 16221 16065 16255 16099
rect 16255 16065 16264 16099
rect 16212 16056 16264 16065
rect 15016 15988 15068 16040
rect 13544 15920 13596 15972
rect 15200 15920 15252 15972
rect 10508 15895 10560 15904
rect 10508 15861 10517 15895
rect 10517 15861 10551 15895
rect 10551 15861 10560 15895
rect 10508 15852 10560 15861
rect 11612 15895 11664 15904
rect 11612 15861 11621 15895
rect 11621 15861 11655 15895
rect 11655 15861 11664 15895
rect 11612 15852 11664 15861
rect 14556 15895 14608 15904
rect 14556 15861 14565 15895
rect 14565 15861 14599 15895
rect 14599 15861 14608 15895
rect 14556 15852 14608 15861
rect 14924 15852 14976 15904
rect 15936 15895 15988 15904
rect 15936 15861 15945 15895
rect 15945 15861 15979 15895
rect 15979 15861 15988 15895
rect 15936 15852 15988 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 4344 15648 4396 15700
rect 4160 15580 4212 15632
rect 1768 15555 1820 15564
rect 1768 15521 1777 15555
rect 1777 15521 1811 15555
rect 1811 15521 1820 15555
rect 1768 15512 1820 15521
rect 2872 15512 2924 15564
rect 4896 15580 4948 15632
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2688 15444 2740 15496
rect 4620 15512 4672 15564
rect 4344 15487 4396 15496
rect 4344 15453 4353 15487
rect 4353 15453 4387 15487
rect 4387 15453 4396 15487
rect 4344 15444 4396 15453
rect 4712 15487 4764 15496
rect 4712 15453 4721 15487
rect 4721 15453 4755 15487
rect 4755 15453 4764 15487
rect 4712 15444 4764 15453
rect 4804 15487 4856 15496
rect 4804 15453 4813 15487
rect 4813 15453 4847 15487
rect 4847 15453 4856 15487
rect 4804 15444 4856 15453
rect 6000 15648 6052 15700
rect 9496 15691 9548 15700
rect 9496 15657 9505 15691
rect 9505 15657 9539 15691
rect 9539 15657 9548 15691
rect 9496 15648 9548 15657
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 17776 15648 17828 15700
rect 11520 15580 11572 15632
rect 12440 15580 12492 15632
rect 12716 15580 12768 15632
rect 6920 15512 6972 15564
rect 10048 15512 10100 15564
rect 10508 15555 10560 15564
rect 10508 15521 10517 15555
rect 10517 15521 10551 15555
rect 10551 15521 10560 15555
rect 10508 15512 10560 15521
rect 4528 15376 4580 15428
rect 6276 15487 6328 15496
rect 6276 15453 6285 15487
rect 6285 15453 6319 15487
rect 6319 15453 6328 15487
rect 6276 15444 6328 15453
rect 6368 15376 6420 15428
rect 7656 15376 7708 15428
rect 9128 15376 9180 15428
rect 9772 15376 9824 15428
rect 11612 15444 11664 15496
rect 12716 15487 12768 15496
rect 12716 15453 12725 15487
rect 12725 15453 12759 15487
rect 12759 15453 12768 15487
rect 12716 15444 12768 15453
rect 13452 15444 13504 15496
rect 16212 15580 16264 15632
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 10416 15376 10468 15428
rect 13176 15376 13228 15428
rect 17316 15444 17368 15496
rect 16580 15376 16632 15428
rect 17960 15376 18012 15428
rect 5356 15308 5408 15360
rect 6092 15351 6144 15360
rect 6092 15317 6101 15351
rect 6101 15317 6135 15351
rect 6135 15317 6144 15351
rect 6092 15308 6144 15317
rect 12900 15308 12952 15360
rect 17592 15351 17644 15360
rect 17592 15317 17601 15351
rect 17601 15317 17635 15351
rect 17635 15317 17644 15351
rect 17592 15308 17644 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 1676 15104 1728 15156
rect 848 14968 900 15020
rect 4344 15104 4396 15156
rect 8576 15104 8628 15156
rect 9036 15147 9088 15156
rect 9036 15113 9045 15147
rect 9045 15113 9079 15147
rect 9079 15113 9088 15147
rect 9036 15104 9088 15113
rect 10048 15104 10100 15156
rect 10876 15147 10928 15156
rect 10876 15113 10885 15147
rect 10885 15113 10919 15147
rect 10919 15113 10928 15147
rect 10876 15104 10928 15113
rect 10968 15104 11020 15156
rect 11244 15104 11296 15156
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 3332 15011 3384 15020
rect 3332 14977 3341 15011
rect 3341 14977 3375 15011
rect 3375 14977 3384 15011
rect 3332 14968 3384 14977
rect 3516 15011 3568 15020
rect 3516 14977 3525 15011
rect 3525 14977 3559 15011
rect 3559 14977 3568 15011
rect 3516 14968 3568 14977
rect 3700 15011 3752 15020
rect 3700 14977 3709 15011
rect 3709 14977 3743 15011
rect 3743 14977 3752 15011
rect 3700 14968 3752 14977
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 4620 15036 4672 15088
rect 5816 15079 5868 15088
rect 5816 15045 5825 15079
rect 5825 15045 5859 15079
rect 5859 15045 5868 15079
rect 5816 15036 5868 15045
rect 6000 15079 6052 15088
rect 6000 15045 6025 15079
rect 6025 15045 6052 15079
rect 6000 15036 6052 15045
rect 4528 15011 4580 15020
rect 4528 14977 4537 15011
rect 4537 14977 4571 15011
rect 4571 14977 4580 15011
rect 4528 14968 4580 14977
rect 6736 15036 6788 15088
rect 7656 15036 7708 15088
rect 11336 15036 11388 15088
rect 1676 14943 1728 14952
rect 1676 14909 1685 14943
rect 1685 14909 1719 14943
rect 1719 14909 1728 14943
rect 1676 14900 1728 14909
rect 1768 14900 1820 14952
rect 2228 14832 2280 14884
rect 3608 14943 3660 14952
rect 3608 14909 3617 14943
rect 3617 14909 3651 14943
rect 3651 14909 3660 14943
rect 3608 14900 3660 14909
rect 4252 14900 4304 14952
rect 3056 14807 3108 14816
rect 3056 14773 3065 14807
rect 3065 14773 3099 14807
rect 3099 14773 3108 14807
rect 3056 14764 3108 14773
rect 4068 14807 4120 14816
rect 4068 14773 4077 14807
rect 4077 14773 4111 14807
rect 4111 14773 4120 14807
rect 4068 14764 4120 14773
rect 4896 14900 4948 14952
rect 5080 14943 5132 14952
rect 5080 14909 5089 14943
rect 5089 14909 5123 14943
rect 5123 14909 5132 14943
rect 5080 14900 5132 14909
rect 4528 14832 4580 14884
rect 5264 14832 5316 14884
rect 4620 14764 4672 14816
rect 4712 14764 4764 14816
rect 6092 14764 6144 14816
rect 6368 14764 6420 14816
rect 9588 15011 9640 15020
rect 9588 14977 9597 15011
rect 9597 14977 9631 15011
rect 9631 14977 9640 15011
rect 9588 14968 9640 14977
rect 11980 15036 12032 15088
rect 12532 14968 12584 15020
rect 13268 15104 13320 15156
rect 13544 15104 13596 15156
rect 15476 15036 15528 15088
rect 9864 14900 9916 14952
rect 11060 14900 11112 14952
rect 11520 14900 11572 14952
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 12440 14900 12492 14952
rect 13544 15011 13596 15020
rect 13544 14977 13553 15011
rect 13553 14977 13587 15011
rect 13587 14977 13596 15011
rect 13544 14968 13596 14977
rect 15384 14968 15436 15020
rect 16672 15011 16724 15020
rect 16672 14977 16681 15011
rect 16681 14977 16715 15011
rect 16715 14977 16724 15011
rect 16672 14968 16724 14977
rect 17040 14968 17092 15020
rect 17408 15036 17460 15088
rect 17592 15147 17644 15156
rect 17592 15113 17601 15147
rect 17601 15113 17635 15147
rect 17635 15113 17644 15147
rect 17592 15104 17644 15113
rect 17776 15104 17828 15156
rect 17224 15011 17276 15020
rect 17224 14977 17233 15011
rect 17233 14977 17267 15011
rect 17267 14977 17276 15011
rect 17224 14968 17276 14977
rect 9956 14832 10008 14884
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 9772 14764 9824 14816
rect 10232 14764 10284 14816
rect 12440 14807 12492 14816
rect 12440 14773 12449 14807
rect 12449 14773 12483 14807
rect 12483 14773 12492 14807
rect 12440 14764 12492 14773
rect 15476 14875 15528 14884
rect 15476 14841 15485 14875
rect 15485 14841 15519 14875
rect 15519 14841 15528 14875
rect 15476 14832 15528 14841
rect 16672 14832 16724 14884
rect 18052 14968 18104 15020
rect 18328 15011 18380 15020
rect 18328 14977 18337 15011
rect 18337 14977 18371 15011
rect 18371 14977 18380 15011
rect 18328 14968 18380 14977
rect 18420 15011 18472 15020
rect 18420 14977 18429 15011
rect 18429 14977 18463 15011
rect 18463 14977 18472 15011
rect 18420 14968 18472 14977
rect 17960 14875 18012 14884
rect 17960 14841 17969 14875
rect 17969 14841 18003 14875
rect 18003 14841 18012 14875
rect 17960 14832 18012 14841
rect 12808 14764 12860 14816
rect 15292 14764 15344 14816
rect 15844 14807 15896 14816
rect 15844 14773 15853 14807
rect 15853 14773 15887 14807
rect 15887 14773 15896 14807
rect 15844 14764 15896 14773
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 2228 14560 2280 14612
rect 2964 14560 3016 14612
rect 3884 14560 3936 14612
rect 3976 14603 4028 14612
rect 3976 14569 3985 14603
rect 3985 14569 4019 14603
rect 4019 14569 4028 14603
rect 3976 14560 4028 14569
rect 4620 14560 4672 14612
rect 4804 14603 4856 14612
rect 4804 14569 4813 14603
rect 4813 14569 4847 14603
rect 4847 14569 4856 14603
rect 4804 14560 4856 14569
rect 5080 14603 5132 14612
rect 5080 14569 5089 14603
rect 5089 14569 5123 14603
rect 5123 14569 5132 14603
rect 5080 14560 5132 14569
rect 6000 14603 6052 14612
rect 6000 14569 6009 14603
rect 6009 14569 6043 14603
rect 6043 14569 6052 14603
rect 6000 14560 6052 14569
rect 1676 14492 1728 14544
rect 2044 14492 2096 14544
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 3056 14424 3108 14476
rect 848 14356 900 14408
rect 3884 14356 3936 14408
rect 5816 14492 5868 14544
rect 6368 14492 6420 14544
rect 6736 14603 6788 14612
rect 6736 14569 6745 14603
rect 6745 14569 6779 14603
rect 6779 14569 6788 14603
rect 6736 14560 6788 14569
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 12440 14560 12492 14612
rect 13452 14560 13504 14612
rect 15476 14560 15528 14612
rect 15752 14560 15804 14612
rect 16672 14603 16724 14612
rect 16672 14569 16681 14603
rect 16681 14569 16715 14603
rect 16715 14569 16724 14603
rect 16672 14560 16724 14569
rect 17224 14560 17276 14612
rect 8668 14492 8720 14544
rect 12532 14492 12584 14544
rect 17408 14560 17460 14612
rect 18328 14560 18380 14612
rect 4620 14424 4672 14476
rect 3608 14288 3660 14340
rect 4804 14356 4856 14408
rect 10876 14424 10928 14476
rect 6276 14356 6328 14408
rect 13268 14424 13320 14476
rect 13360 14424 13412 14476
rect 5448 14288 5500 14340
rect 9588 14288 9640 14340
rect 3976 14220 4028 14272
rect 5816 14220 5868 14272
rect 10324 14331 10376 14340
rect 10324 14297 10333 14331
rect 10333 14297 10367 14331
rect 10367 14297 10376 14331
rect 10324 14288 10376 14297
rect 10416 14263 10468 14272
rect 10416 14229 10425 14263
rect 10425 14229 10459 14263
rect 10459 14229 10468 14263
rect 10416 14220 10468 14229
rect 12808 14288 12860 14340
rect 13452 14356 13504 14408
rect 15936 14467 15988 14476
rect 15936 14433 15945 14467
rect 15945 14433 15979 14467
rect 15979 14433 15988 14467
rect 15936 14424 15988 14433
rect 16396 14467 16448 14476
rect 16396 14433 16405 14467
rect 16405 14433 16439 14467
rect 16439 14433 16448 14467
rect 16396 14424 16448 14433
rect 17960 14492 18012 14544
rect 17776 14424 17828 14476
rect 12072 14220 12124 14272
rect 12992 14263 13044 14272
rect 12992 14229 13001 14263
rect 13001 14229 13035 14263
rect 13035 14229 13044 14263
rect 12992 14220 13044 14229
rect 13728 14331 13780 14340
rect 13728 14297 13737 14331
rect 13737 14297 13771 14331
rect 13771 14297 13780 14331
rect 13728 14288 13780 14297
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 16212 14399 16264 14408
rect 16212 14365 16221 14399
rect 16221 14365 16255 14399
rect 16255 14365 16264 14399
rect 16212 14356 16264 14365
rect 17040 14399 17092 14408
rect 17040 14365 17049 14399
rect 17049 14365 17083 14399
rect 17083 14365 17092 14399
rect 17040 14356 17092 14365
rect 16580 14288 16632 14340
rect 17316 14331 17368 14340
rect 17316 14297 17343 14331
rect 17343 14297 17368 14331
rect 17316 14288 17368 14297
rect 18420 14424 18472 14476
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 17960 14331 18012 14340
rect 17960 14297 17969 14331
rect 17969 14297 18003 14331
rect 18003 14297 18012 14331
rect 17960 14288 18012 14297
rect 16672 14263 16724 14272
rect 16672 14229 16681 14263
rect 16681 14229 16715 14263
rect 16715 14229 16724 14263
rect 16672 14220 16724 14229
rect 17868 14220 17920 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 5816 14059 5868 14068
rect 5816 14025 5825 14059
rect 5825 14025 5859 14059
rect 5859 14025 5868 14059
rect 5816 14016 5868 14025
rect 6368 14016 6420 14068
rect 7656 14016 7708 14068
rect 9864 14016 9916 14068
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 6276 13948 6328 14000
rect 6736 13948 6788 14000
rect 8668 13948 8720 14000
rect 9128 13991 9180 14000
rect 9128 13957 9153 13991
rect 9153 13957 9180 13991
rect 9128 13948 9180 13957
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 2136 13880 2188 13932
rect 2596 13880 2648 13932
rect 5724 13923 5776 13932
rect 5724 13889 5733 13923
rect 5733 13889 5767 13923
rect 5767 13889 5776 13923
rect 5724 13880 5776 13889
rect 6552 13880 6604 13932
rect 7748 13880 7800 13932
rect 10416 13948 10468 14000
rect 12072 13948 12124 14000
rect 16672 14016 16724 14068
rect 16764 14016 16816 14068
rect 18328 14016 18380 14068
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 12624 13948 12676 14000
rect 12992 13948 13044 14000
rect 13176 13948 13228 14000
rect 10508 13812 10560 13864
rect 12072 13812 12124 13864
rect 10692 13744 10744 13796
rect 12440 13812 12492 13864
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 12808 13923 12860 13932
rect 12808 13889 12817 13923
rect 12817 13889 12851 13923
rect 12851 13889 12860 13923
rect 12808 13880 12860 13889
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 13452 13923 13504 13932
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 13452 13880 13504 13889
rect 13084 13744 13136 13796
rect 15108 13923 15160 13932
rect 15108 13889 15117 13923
rect 15117 13889 15151 13923
rect 15151 13889 15160 13923
rect 15108 13880 15160 13889
rect 15200 13880 15252 13932
rect 13820 13855 13872 13864
rect 13820 13821 13829 13855
rect 13829 13821 13863 13855
rect 13863 13821 13872 13855
rect 16120 13880 16172 13932
rect 13820 13812 13872 13821
rect 17040 13812 17092 13864
rect 17868 13880 17920 13932
rect 17776 13855 17828 13864
rect 17776 13821 17785 13855
rect 17785 13821 17819 13855
rect 17819 13821 17828 13855
rect 17776 13812 17828 13821
rect 2596 13676 2648 13728
rect 6368 13676 6420 13728
rect 8668 13676 8720 13728
rect 9220 13676 9272 13728
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 10324 13719 10376 13728
rect 10324 13685 10333 13719
rect 10333 13685 10367 13719
rect 10367 13685 10376 13719
rect 10324 13676 10376 13685
rect 10968 13676 11020 13728
rect 12992 13676 13044 13728
rect 17684 13744 17736 13796
rect 13820 13676 13872 13728
rect 17500 13719 17552 13728
rect 17500 13685 17509 13719
rect 17509 13685 17543 13719
rect 17543 13685 17552 13719
rect 17500 13676 17552 13685
rect 17868 13719 17920 13728
rect 17868 13685 17877 13719
rect 17877 13685 17911 13719
rect 17911 13685 17920 13719
rect 17868 13676 17920 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 4804 13472 4856 13524
rect 5816 13472 5868 13524
rect 6368 13515 6420 13524
rect 6368 13481 6377 13515
rect 6377 13481 6411 13515
rect 6411 13481 6420 13515
rect 6368 13472 6420 13481
rect 6552 13472 6604 13524
rect 8668 13515 8720 13524
rect 8668 13481 8677 13515
rect 8677 13481 8711 13515
rect 8711 13481 8720 13515
rect 8668 13472 8720 13481
rect 10692 13515 10744 13524
rect 2596 13447 2648 13456
rect 2596 13413 2605 13447
rect 2605 13413 2639 13447
rect 2639 13413 2648 13447
rect 2596 13404 2648 13413
rect 3332 13404 3384 13456
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 2044 13336 2096 13388
rect 2688 13336 2740 13388
rect 2136 13311 2188 13320
rect 2136 13277 2145 13311
rect 2145 13277 2179 13311
rect 2179 13277 2188 13311
rect 2136 13268 2188 13277
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 3976 13336 4028 13388
rect 3516 13268 3568 13320
rect 3884 13311 3936 13320
rect 3884 13277 3893 13311
rect 3893 13277 3927 13311
rect 3927 13277 3936 13311
rect 3884 13268 3936 13277
rect 3240 13243 3292 13252
rect 3240 13209 3249 13243
rect 3249 13209 3283 13243
rect 3283 13209 3292 13243
rect 3240 13200 3292 13209
rect 6644 13379 6696 13388
rect 6644 13345 6653 13379
rect 6653 13345 6687 13379
rect 6687 13345 6696 13379
rect 6644 13336 6696 13345
rect 4160 13243 4212 13252
rect 4160 13209 4169 13243
rect 4169 13209 4203 13243
rect 4203 13209 4212 13243
rect 4160 13200 4212 13209
rect 5632 13200 5684 13252
rect 5724 13243 5776 13252
rect 5724 13209 5749 13243
rect 5749 13209 5776 13243
rect 5724 13200 5776 13209
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 12808 13472 12860 13524
rect 12716 13404 12768 13456
rect 10876 13379 10928 13388
rect 10876 13345 10885 13379
rect 10885 13345 10919 13379
rect 10919 13345 10928 13379
rect 10876 13336 10928 13345
rect 848 13132 900 13184
rect 2228 13132 2280 13184
rect 3976 13132 4028 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 7932 13200 7984 13252
rect 12624 13268 12676 13320
rect 12992 13311 13044 13320
rect 12992 13277 13001 13311
rect 13001 13277 13035 13311
rect 13035 13277 13044 13311
rect 12992 13268 13044 13277
rect 13728 13515 13780 13524
rect 13728 13481 13737 13515
rect 13737 13481 13771 13515
rect 13771 13481 13780 13515
rect 13728 13472 13780 13481
rect 17316 13472 17368 13524
rect 16580 13336 16632 13388
rect 17684 13336 17736 13388
rect 9220 13243 9272 13252
rect 9220 13209 9229 13243
rect 9229 13209 9263 13243
rect 9263 13209 9272 13243
rect 9220 13200 9272 13209
rect 9772 13200 9824 13252
rect 11152 13243 11204 13252
rect 11152 13209 11161 13243
rect 11161 13209 11195 13243
rect 11195 13209 11204 13243
rect 11152 13200 11204 13209
rect 11796 13200 11848 13252
rect 13084 13200 13136 13252
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 13820 13311 13872 13320
rect 13820 13277 13829 13311
rect 13829 13277 13863 13311
rect 13863 13277 13872 13311
rect 13820 13268 13872 13277
rect 17500 13268 17552 13320
rect 18512 13311 18564 13320
rect 18512 13277 18521 13311
rect 18521 13277 18555 13311
rect 18555 13277 18564 13311
rect 18512 13268 18564 13277
rect 15200 13200 15252 13252
rect 9864 13132 9916 13184
rect 12072 13132 12124 13184
rect 13728 13132 13780 13184
rect 18420 13132 18472 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 3240 12928 3292 12980
rect 2044 12835 2096 12844
rect 2044 12801 2053 12835
rect 2053 12801 2087 12835
rect 2087 12801 2096 12835
rect 2044 12792 2096 12801
rect 2228 12724 2280 12776
rect 1584 12656 1636 12708
rect 2688 12724 2740 12776
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 5632 12971 5684 12980
rect 5632 12937 5641 12971
rect 5641 12937 5675 12971
rect 5675 12937 5684 12971
rect 5632 12928 5684 12937
rect 5724 12928 5776 12980
rect 5908 12928 5960 12980
rect 2964 12724 3016 12776
rect 3884 12724 3936 12776
rect 4712 12792 4764 12844
rect 6368 12860 6420 12912
rect 7932 12928 7984 12980
rect 9128 12928 9180 12980
rect 9680 12928 9732 12980
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 11152 12928 11204 12980
rect 11796 12971 11848 12980
rect 11796 12937 11805 12971
rect 11805 12937 11839 12971
rect 11839 12937 11848 12971
rect 11796 12928 11848 12937
rect 12440 12928 12492 12980
rect 13544 12928 13596 12980
rect 15660 12928 15712 12980
rect 16120 12971 16172 12980
rect 16120 12937 16129 12971
rect 16129 12937 16163 12971
rect 16163 12937 16172 12971
rect 16120 12928 16172 12937
rect 16580 12928 16632 12980
rect 4620 12724 4672 12776
rect 5540 12792 5592 12844
rect 5816 12792 5868 12844
rect 9864 12860 9916 12912
rect 10692 12903 10744 12912
rect 10692 12869 10701 12903
rect 10701 12869 10735 12903
rect 10735 12869 10744 12903
rect 10692 12860 10744 12869
rect 14004 12860 14056 12912
rect 15016 12860 15068 12912
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7748 12792 7800 12844
rect 7932 12835 7984 12844
rect 7932 12801 7941 12835
rect 7941 12801 7975 12835
rect 7975 12801 7984 12835
rect 7932 12792 7984 12801
rect 3056 12656 3108 12708
rect 3976 12656 4028 12708
rect 4068 12656 4120 12708
rect 4988 12767 5040 12776
rect 4988 12733 4997 12767
rect 4997 12733 5031 12767
rect 5031 12733 5040 12767
rect 4988 12724 5040 12733
rect 10140 12724 10192 12776
rect 10324 12835 10376 12844
rect 10324 12801 10333 12835
rect 10333 12801 10367 12835
rect 10367 12801 10376 12835
rect 10324 12792 10376 12801
rect 11060 12724 11112 12776
rect 13360 12792 13412 12844
rect 17500 12860 17552 12912
rect 13820 12724 13872 12776
rect 1676 12631 1728 12640
rect 1676 12597 1685 12631
rect 1685 12597 1719 12631
rect 1719 12597 1728 12631
rect 1676 12588 1728 12597
rect 2136 12588 2188 12640
rect 2872 12588 2924 12640
rect 5908 12588 5960 12640
rect 14648 12656 14700 12708
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 16120 12724 16172 12776
rect 16580 12724 16632 12776
rect 16764 12792 16816 12844
rect 17408 12835 17460 12844
rect 17408 12801 17417 12835
rect 17417 12801 17451 12835
rect 17451 12801 17460 12835
rect 17408 12792 17460 12801
rect 18420 12835 18472 12844
rect 16028 12656 16080 12708
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 18420 12801 18429 12835
rect 18429 12801 18463 12835
rect 18463 12801 18472 12835
rect 18420 12792 18472 12801
rect 6920 12631 6972 12640
rect 6920 12597 6929 12631
rect 6929 12597 6963 12631
rect 6963 12597 6972 12631
rect 6920 12588 6972 12597
rect 11980 12588 12032 12640
rect 14740 12588 14792 12640
rect 15200 12588 15252 12640
rect 15660 12588 15712 12640
rect 17592 12631 17644 12640
rect 17592 12597 17616 12631
rect 17616 12597 17644 12631
rect 17592 12588 17644 12597
rect 17684 12631 17736 12640
rect 17684 12597 17693 12631
rect 17693 12597 17727 12631
rect 17727 12597 17736 12631
rect 17684 12588 17736 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 3792 12384 3844 12436
rect 2504 12316 2556 12368
rect 3424 12316 3476 12368
rect 1676 12248 1728 12300
rect 4160 12291 4212 12300
rect 848 12180 900 12232
rect 2228 12180 2280 12232
rect 2596 12180 2648 12232
rect 2504 12112 2556 12164
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 4160 12257 4169 12291
rect 4169 12257 4203 12291
rect 4203 12257 4212 12291
rect 4160 12248 4212 12257
rect 3976 12180 4028 12232
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4712 12223 4764 12232
rect 4436 12180 4488 12189
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 4988 12180 5040 12232
rect 5356 12384 5408 12436
rect 7196 12384 7248 12436
rect 10692 12384 10744 12436
rect 14464 12427 14516 12436
rect 14464 12393 14473 12427
rect 14473 12393 14507 12427
rect 14507 12393 14516 12427
rect 14464 12384 14516 12393
rect 5356 12248 5408 12300
rect 7932 12248 7984 12300
rect 2964 12044 3016 12096
rect 3976 12044 4028 12096
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 6460 12180 6512 12189
rect 9680 12248 9732 12300
rect 14648 12291 14700 12300
rect 14648 12257 14657 12291
rect 14657 12257 14691 12291
rect 14691 12257 14700 12291
rect 14648 12248 14700 12257
rect 15936 12384 15988 12436
rect 16120 12427 16172 12436
rect 16120 12393 16129 12427
rect 16129 12393 16163 12427
rect 16163 12393 16172 12427
rect 16120 12384 16172 12393
rect 17040 12384 17092 12436
rect 15108 12359 15160 12368
rect 15108 12325 15117 12359
rect 15117 12325 15151 12359
rect 15151 12325 15160 12359
rect 15108 12316 15160 12325
rect 15200 12248 15252 12300
rect 9864 12180 9916 12232
rect 10140 12223 10192 12232
rect 10140 12189 10149 12223
rect 10149 12189 10183 12223
rect 10183 12189 10192 12223
rect 10140 12180 10192 12189
rect 10508 12180 10560 12232
rect 11336 12180 11388 12232
rect 5264 12044 5316 12096
rect 5448 12087 5500 12096
rect 5448 12053 5457 12087
rect 5457 12053 5491 12087
rect 5491 12053 5500 12087
rect 5448 12044 5500 12053
rect 6920 12044 6972 12096
rect 11888 12087 11940 12096
rect 11888 12053 11897 12087
rect 11897 12053 11931 12087
rect 11931 12053 11940 12087
rect 11888 12044 11940 12053
rect 15016 12180 15068 12232
rect 15660 12248 15712 12300
rect 15936 12223 15988 12232
rect 15936 12189 15945 12223
rect 15945 12189 15979 12223
rect 15979 12189 15988 12223
rect 15936 12180 15988 12189
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 17408 12180 17460 12232
rect 17684 12180 17736 12232
rect 18512 12223 18564 12232
rect 18512 12189 18521 12223
rect 18521 12189 18555 12223
rect 18555 12189 18564 12223
rect 18512 12180 18564 12189
rect 16764 12112 16816 12164
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2044 11840 2096 11892
rect 2688 11840 2740 11892
rect 4436 11840 4488 11892
rect 5448 11840 5500 11892
rect 848 11704 900 11756
rect 7932 11772 7984 11824
rect 8024 11815 8076 11824
rect 8024 11781 8033 11815
rect 8033 11781 8067 11815
rect 8067 11781 8076 11815
rect 8024 11772 8076 11781
rect 9588 11815 9640 11824
rect 9588 11781 9597 11815
rect 9597 11781 9631 11815
rect 9631 11781 9640 11815
rect 9588 11772 9640 11781
rect 12532 11840 12584 11892
rect 11796 11772 11848 11824
rect 11888 11772 11940 11824
rect 1584 11636 1636 11688
rect 4068 11747 4120 11756
rect 4068 11713 4078 11747
rect 4078 11713 4112 11747
rect 4112 11713 4120 11747
rect 4068 11704 4120 11713
rect 9864 11747 9916 11756
rect 9864 11713 9873 11747
rect 9873 11713 9907 11747
rect 9907 11713 9916 11747
rect 9864 11704 9916 11713
rect 10140 11704 10192 11756
rect 10876 11704 10928 11756
rect 4620 11636 4672 11688
rect 9956 11636 10008 11688
rect 10784 11636 10836 11688
rect 2136 11543 2188 11552
rect 2136 11509 2145 11543
rect 2145 11509 2179 11543
rect 2179 11509 2188 11543
rect 2136 11500 2188 11509
rect 5540 11500 5592 11552
rect 9128 11568 9180 11620
rect 13268 11636 13320 11688
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14096 11747 14148 11756
rect 14096 11713 14105 11747
rect 14105 11713 14139 11747
rect 14139 11713 14148 11747
rect 14096 11704 14148 11713
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16856 11704 16908 11756
rect 16948 11636 17000 11688
rect 8944 11500 8996 11552
rect 9312 11500 9364 11552
rect 10232 11500 10284 11552
rect 13544 11500 13596 11552
rect 13820 11543 13872 11552
rect 13820 11509 13829 11543
rect 13829 11509 13863 11543
rect 13863 11509 13872 11543
rect 13820 11500 13872 11509
rect 13912 11500 13964 11552
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 16028 11500 16080 11552
rect 16764 11500 16816 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 5356 11296 5408 11348
rect 5540 11339 5592 11348
rect 5540 11305 5549 11339
rect 5549 11305 5583 11339
rect 5583 11305 5592 11339
rect 5540 11296 5592 11305
rect 10784 11339 10836 11348
rect 10784 11305 10793 11339
rect 10793 11305 10827 11339
rect 10827 11305 10836 11339
rect 10784 11296 10836 11305
rect 11796 11339 11848 11348
rect 11796 11305 11805 11339
rect 11805 11305 11839 11339
rect 11839 11305 11848 11339
rect 11796 11296 11848 11305
rect 14096 11296 14148 11348
rect 15752 11296 15804 11348
rect 8576 11228 8628 11280
rect 6460 11160 6512 11212
rect 6552 11160 6604 11212
rect 9312 11203 9364 11212
rect 9312 11169 9321 11203
rect 9321 11169 9355 11203
rect 9355 11169 9364 11203
rect 9312 11160 9364 11169
rect 3424 11092 3476 11144
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 4252 11092 4304 11144
rect 4436 11135 4488 11144
rect 4436 11101 4445 11135
rect 4445 11101 4479 11135
rect 4479 11101 4488 11135
rect 4436 11092 4488 11101
rect 4620 11135 4672 11144
rect 4620 11101 4633 11135
rect 4633 11101 4672 11135
rect 4620 11092 4672 11101
rect 5356 11092 5408 11144
rect 7932 11135 7984 11144
rect 7932 11101 7941 11135
rect 7941 11101 7975 11135
rect 7975 11101 7984 11135
rect 7932 11092 7984 11101
rect 9128 11135 9180 11144
rect 9128 11101 9137 11135
rect 9137 11101 9171 11135
rect 9171 11101 9180 11135
rect 9128 11092 9180 11101
rect 12900 11228 12952 11280
rect 13912 11160 13964 11212
rect 16304 11228 16356 11280
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 10048 11135 10100 11144
rect 10048 11101 10057 11135
rect 10057 11101 10091 11135
rect 10091 11101 10100 11135
rect 10048 11092 10100 11101
rect 2136 11024 2188 11076
rect 4068 11067 4120 11076
rect 4068 11033 4077 11067
rect 4077 11033 4111 11067
rect 4111 11033 4120 11067
rect 4068 11024 4120 11033
rect 5632 11024 5684 11076
rect 4160 10956 4212 11008
rect 8668 11024 8720 11076
rect 9404 11024 9456 11076
rect 10968 11092 11020 11144
rect 11244 11024 11296 11076
rect 11428 11067 11480 11076
rect 11428 11033 11437 11067
rect 11437 11033 11471 11067
rect 11471 11033 11480 11067
rect 11428 11024 11480 11033
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 13360 11135 13412 11144
rect 13360 11101 13369 11135
rect 13369 11101 13403 11135
rect 13403 11101 13412 11135
rect 13360 11092 13412 11101
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 14004 11092 14056 11144
rect 15292 11092 15344 11144
rect 15844 11092 15896 11144
rect 10692 10956 10744 11008
rect 11152 10999 11204 11008
rect 11152 10965 11161 10999
rect 11161 10965 11195 10999
rect 11195 10965 11204 10999
rect 11152 10956 11204 10965
rect 12348 10956 12400 11008
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 16396 11024 16448 11076
rect 16120 10956 16172 11008
rect 16856 11024 16908 11076
rect 16948 11067 17000 11076
rect 16948 11033 16957 11067
rect 16957 11033 16991 11067
rect 16991 11033 17000 11067
rect 16948 11024 17000 11033
rect 17224 10956 17276 11008
rect 17960 10956 18012 11008
rect 18236 11135 18288 11144
rect 18236 11101 18245 11135
rect 18245 11101 18279 11135
rect 18279 11101 18288 11135
rect 18236 11092 18288 11101
rect 18512 11135 18564 11144
rect 18512 11101 18521 11135
rect 18521 11101 18555 11135
rect 18555 11101 18564 11135
rect 18512 11092 18564 11101
rect 18328 10999 18380 11008
rect 18328 10965 18337 10999
rect 18337 10965 18371 10999
rect 18371 10965 18380 10999
rect 18328 10956 18380 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 4252 10752 4304 10804
rect 5540 10795 5592 10804
rect 5540 10761 5549 10795
rect 5549 10761 5583 10795
rect 5583 10761 5592 10795
rect 5540 10752 5592 10761
rect 10048 10752 10100 10804
rect 848 10616 900 10668
rect 2688 10616 2740 10668
rect 4712 10684 4764 10736
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 4804 10616 4856 10668
rect 5448 10684 5500 10736
rect 5908 10727 5960 10736
rect 5908 10693 5917 10727
rect 5917 10693 5951 10727
rect 5951 10693 5960 10727
rect 5908 10684 5960 10693
rect 6552 10684 6604 10736
rect 9680 10727 9732 10736
rect 9680 10693 9689 10727
rect 9689 10693 9723 10727
rect 9723 10693 9732 10727
rect 9680 10684 9732 10693
rect 2596 10548 2648 10600
rect 3884 10548 3936 10600
rect 4528 10548 4580 10600
rect 7748 10616 7800 10668
rect 5264 10412 5316 10464
rect 5356 10412 5408 10464
rect 6644 10591 6696 10600
rect 6644 10557 6653 10591
rect 6653 10557 6687 10591
rect 6687 10557 6696 10591
rect 6644 10548 6696 10557
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 11428 10752 11480 10804
rect 13176 10752 13228 10804
rect 13452 10752 13504 10804
rect 14648 10752 14700 10804
rect 10140 10548 10192 10600
rect 10692 10659 10744 10668
rect 10692 10625 10701 10659
rect 10701 10625 10735 10659
rect 10735 10625 10744 10659
rect 10692 10616 10744 10625
rect 10876 10684 10928 10736
rect 11152 10616 11204 10668
rect 15016 10684 15068 10736
rect 12348 10659 12400 10668
rect 12348 10625 12357 10659
rect 12357 10625 12391 10659
rect 12391 10625 12400 10659
rect 12348 10616 12400 10625
rect 13176 10616 13228 10668
rect 8852 10523 8904 10532
rect 8852 10489 8861 10523
rect 8861 10489 8895 10523
rect 8895 10489 8904 10523
rect 8852 10480 8904 10489
rect 13820 10548 13872 10600
rect 7104 10412 7156 10464
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 9496 10455 9548 10464
rect 9496 10421 9505 10455
rect 9505 10421 9539 10455
rect 9539 10421 9548 10455
rect 9496 10412 9548 10421
rect 10968 10455 11020 10464
rect 10968 10421 10977 10455
rect 10977 10421 11011 10455
rect 11011 10421 11020 10455
rect 10968 10412 11020 10421
rect 13084 10455 13136 10464
rect 13084 10421 13093 10455
rect 13093 10421 13127 10455
rect 13127 10421 13136 10455
rect 13084 10412 13136 10421
rect 13360 10412 13412 10464
rect 13636 10412 13688 10464
rect 14004 10659 14056 10668
rect 14004 10625 14013 10659
rect 14013 10625 14047 10659
rect 14047 10625 14056 10659
rect 14004 10616 14056 10625
rect 14648 10616 14700 10668
rect 15200 10684 15252 10736
rect 15936 10684 15988 10736
rect 16304 10727 16356 10736
rect 16304 10693 16313 10727
rect 16313 10693 16347 10727
rect 16347 10693 16356 10727
rect 16304 10684 16356 10693
rect 16488 10684 16540 10736
rect 16856 10795 16908 10804
rect 16856 10761 16865 10795
rect 16865 10761 16899 10795
rect 16899 10761 16908 10795
rect 16856 10752 16908 10761
rect 17224 10684 17276 10736
rect 17316 10684 17368 10736
rect 15384 10616 15436 10668
rect 15660 10616 15712 10668
rect 16120 10659 16172 10668
rect 16120 10625 16129 10659
rect 16129 10625 16163 10659
rect 16163 10625 16172 10659
rect 16120 10616 16172 10625
rect 16396 10659 16448 10668
rect 16396 10625 16405 10659
rect 16405 10625 16439 10659
rect 16439 10625 16448 10659
rect 16396 10616 16448 10625
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17224 10591 17276 10600
rect 17224 10557 17233 10591
rect 17233 10557 17267 10591
rect 17267 10557 17276 10591
rect 17224 10548 17276 10557
rect 17592 10548 17644 10600
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 15384 10480 15436 10532
rect 15660 10480 15712 10532
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 16304 10412 16356 10464
rect 17132 10412 17184 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 2688 10251 2740 10260
rect 2688 10217 2697 10251
rect 2697 10217 2731 10251
rect 2731 10217 2740 10251
rect 2688 10208 2740 10217
rect 1860 10072 1912 10124
rect 2596 10072 2648 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 1952 10004 2004 10056
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5356 10208 5408 10260
rect 6092 10004 6144 10056
rect 1676 9868 1728 9920
rect 4620 9868 4672 9920
rect 6000 9868 6052 9920
rect 7748 10208 7800 10260
rect 9496 10208 9548 10260
rect 10140 10208 10192 10260
rect 11152 10208 11204 10260
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 15476 10208 15528 10260
rect 16212 10251 16264 10260
rect 16212 10217 16221 10251
rect 16221 10217 16255 10251
rect 16255 10217 16264 10251
rect 16212 10208 16264 10217
rect 16304 10251 16356 10260
rect 16304 10217 16313 10251
rect 16313 10217 16347 10251
rect 16347 10217 16356 10251
rect 16304 10208 16356 10217
rect 16396 10208 16448 10260
rect 18328 10208 18380 10260
rect 9772 10072 9824 10124
rect 13084 10140 13136 10192
rect 8116 10004 8168 10056
rect 8668 10047 8720 10056
rect 8668 10013 8677 10047
rect 8677 10013 8711 10047
rect 8711 10013 8720 10047
rect 8668 10004 8720 10013
rect 7380 9936 7432 9988
rect 8576 9936 8628 9988
rect 11244 10004 11296 10056
rect 12992 10047 13044 10056
rect 12992 10013 13001 10047
rect 13001 10013 13035 10047
rect 13035 10013 13044 10047
rect 12992 10004 13044 10013
rect 16488 10140 16540 10192
rect 17592 10140 17644 10192
rect 13268 10004 13320 10056
rect 14188 10004 14240 10056
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 15108 10115 15160 10124
rect 15108 10081 15117 10115
rect 15117 10081 15151 10115
rect 15151 10081 15160 10115
rect 15108 10072 15160 10081
rect 15292 10115 15344 10124
rect 15292 10081 15338 10115
rect 15338 10081 15344 10115
rect 15292 10072 15344 10081
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 15200 10004 15252 10056
rect 15752 10047 15804 10056
rect 15752 10013 15761 10047
rect 15761 10013 15795 10047
rect 15795 10013 15804 10047
rect 15752 10004 15804 10013
rect 15384 9936 15436 9988
rect 15936 10047 15988 10056
rect 15936 10013 15945 10047
rect 15945 10013 15979 10047
rect 15979 10013 15988 10047
rect 15936 10004 15988 10013
rect 17960 10072 18012 10124
rect 16396 10047 16448 10056
rect 16396 10013 16405 10047
rect 16405 10013 16439 10047
rect 16439 10013 16448 10047
rect 16396 10004 16448 10013
rect 17224 10004 17276 10056
rect 17316 10047 17368 10056
rect 17316 10013 17325 10047
rect 17325 10013 17359 10047
rect 17359 10013 17368 10047
rect 17316 10004 17368 10013
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 7012 9911 7064 9920
rect 7012 9877 7021 9911
rect 7021 9877 7055 9911
rect 7055 9877 7064 9911
rect 7012 9868 7064 9877
rect 14372 9868 14424 9920
rect 15108 9868 15160 9920
rect 15200 9868 15252 9920
rect 16028 9868 16080 9920
rect 16396 9868 16448 9920
rect 17132 9868 17184 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 1952 9664 2004 9716
rect 6644 9664 6696 9716
rect 1676 9528 1728 9580
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 1584 9392 1636 9444
rect 2964 9460 3016 9512
rect 2228 9435 2280 9444
rect 2228 9401 2237 9435
rect 2237 9401 2271 9435
rect 2271 9401 2280 9435
rect 2228 9392 2280 9401
rect 2320 9324 2372 9376
rect 3148 9324 3200 9376
rect 4068 9528 4120 9580
rect 4712 9596 4764 9648
rect 5632 9596 5684 9648
rect 7012 9596 7064 9648
rect 9680 9596 9732 9648
rect 10416 9639 10468 9648
rect 10416 9605 10425 9639
rect 10425 9605 10459 9639
rect 10459 9605 10468 9639
rect 10416 9596 10468 9605
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10968 9528 11020 9580
rect 12256 9596 12308 9648
rect 13636 9707 13688 9716
rect 13636 9673 13645 9707
rect 13645 9673 13679 9707
rect 13679 9673 13688 9707
rect 13636 9664 13688 9673
rect 13912 9664 13964 9716
rect 14648 9664 14700 9716
rect 15292 9664 15344 9716
rect 15752 9664 15804 9716
rect 18328 9707 18380 9716
rect 18328 9673 18337 9707
rect 18337 9673 18371 9707
rect 18371 9673 18380 9707
rect 18328 9664 18380 9673
rect 15568 9639 15620 9648
rect 11152 9528 11204 9580
rect 15568 9605 15577 9639
rect 15577 9605 15611 9639
rect 15611 9605 15620 9639
rect 15568 9596 15620 9605
rect 17224 9596 17276 9648
rect 13912 9571 13964 9580
rect 13912 9537 13921 9571
rect 13921 9537 13955 9571
rect 13955 9537 13964 9571
rect 13912 9528 13964 9537
rect 3884 9503 3936 9512
rect 3884 9469 3893 9503
rect 3893 9469 3927 9503
rect 3927 9469 3936 9503
rect 3884 9460 3936 9469
rect 9772 9460 9824 9512
rect 3976 9324 4028 9376
rect 4712 9324 4764 9376
rect 6000 9367 6052 9376
rect 6000 9333 6009 9367
rect 6009 9333 6043 9367
rect 6043 9333 6052 9367
rect 6000 9324 6052 9333
rect 14372 9528 14424 9580
rect 14280 9460 14332 9512
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 15660 9571 15712 9580
rect 15660 9537 15674 9571
rect 15674 9537 15708 9571
rect 15708 9537 15712 9571
rect 15660 9528 15712 9537
rect 17960 9571 18012 9580
rect 17960 9537 17969 9571
rect 17969 9537 18003 9571
rect 18003 9537 18012 9571
rect 17960 9528 18012 9537
rect 18512 9571 18564 9580
rect 18512 9537 18521 9571
rect 18521 9537 18555 9571
rect 18555 9537 18564 9571
rect 18512 9528 18564 9537
rect 16028 9460 16080 9512
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 13820 9392 13872 9444
rect 15476 9392 15528 9444
rect 17408 9392 17460 9444
rect 16304 9324 16356 9376
rect 18236 9367 18288 9376
rect 18236 9333 18245 9367
rect 18245 9333 18279 9367
rect 18279 9333 18288 9367
rect 18236 9324 18288 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 848 8916 900 8968
rect 3332 9120 3384 9172
rect 3884 9120 3936 9172
rect 2964 9052 3016 9104
rect 2228 9027 2280 9036
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 2320 8984 2372 9036
rect 5448 9120 5500 9172
rect 8852 9120 8904 9172
rect 10140 9120 10192 9172
rect 10692 9120 10744 9172
rect 10968 9120 11020 9172
rect 12256 9120 12308 9172
rect 15476 9120 15528 9172
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 2780 8916 2832 8925
rect 3516 8984 3568 9036
rect 4620 8984 4672 9036
rect 5080 9052 5132 9104
rect 4896 8984 4948 9036
rect 3056 8891 3108 8900
rect 3056 8857 3065 8891
rect 3065 8857 3099 8891
rect 3099 8857 3108 8891
rect 3056 8848 3108 8857
rect 3148 8848 3200 8900
rect 3792 8916 3844 8968
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4344 8916 4396 8968
rect 4804 8916 4856 8968
rect 2596 8823 2648 8832
rect 2596 8789 2605 8823
rect 2605 8789 2639 8823
rect 2639 8789 2648 8823
rect 2596 8780 2648 8789
rect 3976 8780 4028 8832
rect 5080 8891 5132 8900
rect 5080 8857 5089 8891
rect 5089 8857 5123 8891
rect 5123 8857 5132 8891
rect 5080 8848 5132 8857
rect 6092 8916 6144 8968
rect 6184 8959 6236 8968
rect 6184 8925 6193 8959
rect 6193 8925 6227 8959
rect 6227 8925 6236 8959
rect 6184 8916 6236 8925
rect 8024 8984 8076 9036
rect 8392 9027 8444 9036
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 9128 9052 9180 9104
rect 9036 8984 9088 9036
rect 9496 8984 9548 9036
rect 10600 8984 10652 9036
rect 5448 8891 5500 8900
rect 5448 8857 5457 8891
rect 5457 8857 5491 8891
rect 5491 8857 5500 8891
rect 5448 8848 5500 8857
rect 6276 8848 6328 8900
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 7288 8848 7340 8900
rect 5356 8780 5408 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 7196 8780 7248 8832
rect 8300 8916 8352 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 9220 8848 9272 8900
rect 10140 8848 10192 8900
rect 11244 8916 11296 8968
rect 12164 8916 12216 8968
rect 16856 8916 16908 8968
rect 17316 9120 17368 9172
rect 18052 9120 18104 9172
rect 18512 9120 18564 9172
rect 17224 9027 17276 9036
rect 17224 8993 17233 9027
rect 17233 8993 17267 9027
rect 17267 8993 17276 9027
rect 17224 8984 17276 8993
rect 17408 8916 17460 8968
rect 18328 8984 18380 9036
rect 18236 8959 18288 8968
rect 18236 8925 18245 8959
rect 18245 8925 18279 8959
rect 18279 8925 18288 8959
rect 18236 8916 18288 8925
rect 11336 8848 11388 8900
rect 13544 8848 13596 8900
rect 17684 8891 17736 8900
rect 17684 8857 17718 8891
rect 17718 8857 17736 8891
rect 17684 8848 17736 8857
rect 18052 8848 18104 8900
rect 9864 8780 9916 8832
rect 10784 8780 10836 8832
rect 16212 8780 16264 8832
rect 17224 8780 17276 8832
rect 17592 8823 17644 8832
rect 17592 8789 17601 8823
rect 17601 8789 17635 8823
rect 17635 8789 17644 8823
rect 17592 8780 17644 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2320 8576 2372 8628
rect 1860 8440 1912 8492
rect 3056 8508 3108 8560
rect 2504 8440 2556 8492
rect 4344 8619 4396 8628
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 3608 8508 3660 8560
rect 4896 8576 4948 8628
rect 5172 8576 5224 8628
rect 8300 8619 8352 8628
rect 8300 8585 8309 8619
rect 8309 8585 8343 8619
rect 8343 8585 8352 8619
rect 8300 8576 8352 8585
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 6092 8508 6144 8560
rect 1400 8415 1452 8424
rect 1400 8381 1409 8415
rect 1409 8381 1443 8415
rect 1443 8381 1452 8415
rect 1400 8372 1452 8381
rect 2780 8372 2832 8424
rect 3240 8304 3292 8356
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 5264 8440 5316 8492
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 5632 8372 5684 8424
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6184 8440 6236 8492
rect 6460 8483 6512 8492
rect 6460 8449 6469 8483
rect 6469 8449 6503 8483
rect 6503 8449 6512 8483
rect 6460 8440 6512 8449
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 8024 8508 8076 8560
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7840 8440 7892 8492
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 8484 8440 8536 8492
rect 4712 8304 4764 8356
rect 4896 8304 4948 8356
rect 5448 8304 5500 8356
rect 6460 8304 6512 8356
rect 7196 8372 7248 8424
rect 8208 8372 8260 8424
rect 9404 8576 9456 8628
rect 9496 8576 9548 8628
rect 12992 8576 13044 8628
rect 14004 8576 14056 8628
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 17684 8576 17736 8628
rect 9772 8508 9824 8560
rect 11520 8508 11572 8560
rect 9220 8483 9272 8492
rect 9220 8449 9229 8483
rect 9229 8449 9263 8483
rect 9263 8449 9272 8483
rect 9220 8440 9272 8449
rect 9404 8440 9456 8492
rect 8944 8304 8996 8356
rect 9864 8483 9916 8492
rect 9864 8449 9873 8483
rect 9873 8449 9907 8483
rect 9907 8449 9916 8483
rect 9864 8440 9916 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 14096 8508 14148 8560
rect 18512 8576 18564 8628
rect 9956 8372 10008 8424
rect 10048 8372 10100 8424
rect 10324 8372 10376 8424
rect 13268 8372 13320 8424
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 13912 8483 13964 8492
rect 13912 8449 13921 8483
rect 13921 8449 13955 8483
rect 13955 8449 13964 8483
rect 13912 8440 13964 8449
rect 14372 8440 14424 8492
rect 15476 8440 15528 8492
rect 17040 8440 17092 8492
rect 17500 8440 17552 8492
rect 18420 8551 18472 8560
rect 18420 8517 18429 8551
rect 18429 8517 18463 8551
rect 18463 8517 18472 8551
rect 18420 8508 18472 8517
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 18052 8440 18104 8492
rect 12348 8304 12400 8356
rect 13820 8304 13872 8356
rect 18236 8372 18288 8424
rect 17316 8304 17368 8356
rect 17960 8304 18012 8356
rect 2688 8236 2740 8288
rect 2964 8279 3016 8288
rect 2964 8245 2973 8279
rect 2973 8245 3007 8279
rect 3007 8245 3016 8279
rect 2964 8236 3016 8245
rect 3332 8279 3384 8288
rect 3332 8245 3341 8279
rect 3341 8245 3375 8279
rect 3375 8245 3384 8279
rect 3332 8236 3384 8245
rect 5816 8279 5868 8288
rect 5816 8245 5825 8279
rect 5825 8245 5859 8279
rect 5859 8245 5868 8279
rect 5816 8236 5868 8245
rect 9220 8236 9272 8288
rect 9680 8236 9732 8288
rect 11612 8279 11664 8288
rect 11612 8245 11621 8279
rect 11621 8245 11655 8279
rect 11655 8245 11664 8279
rect 11612 8236 11664 8245
rect 17408 8279 17460 8288
rect 17408 8245 17417 8279
rect 17417 8245 17451 8279
rect 17451 8245 17460 8279
rect 17408 8236 17460 8245
rect 17868 8236 17920 8288
rect 18236 8236 18288 8288
rect 18420 8236 18472 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4068 8032 4120 8084
rect 4620 8032 4672 8084
rect 7932 8032 7984 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 9312 8032 9364 8084
rect 10140 8075 10192 8084
rect 10140 8041 10149 8075
rect 10149 8041 10183 8075
rect 10183 8041 10192 8075
rect 10140 8032 10192 8041
rect 11612 8032 11664 8084
rect 14188 8075 14240 8084
rect 14188 8041 14197 8075
rect 14197 8041 14231 8075
rect 14231 8041 14240 8075
rect 14188 8032 14240 8041
rect 2596 7939 2648 7948
rect 2596 7905 2605 7939
rect 2605 7905 2639 7939
rect 2639 7905 2648 7939
rect 2596 7896 2648 7905
rect 2964 7896 3016 7948
rect 848 7828 900 7880
rect 2504 7871 2556 7880
rect 2504 7837 2513 7871
rect 2513 7837 2547 7871
rect 2547 7837 2556 7871
rect 2504 7828 2556 7837
rect 3240 7828 3292 7880
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4712 7896 4764 7948
rect 2688 7760 2740 7812
rect 4252 7803 4304 7812
rect 4252 7769 4261 7803
rect 4261 7769 4295 7803
rect 4295 7769 4304 7803
rect 4252 7760 4304 7769
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 6828 7964 6880 8016
rect 8208 7964 8260 8016
rect 13912 7964 13964 8016
rect 15108 8007 15160 8016
rect 15108 7973 15117 8007
rect 15117 7973 15151 8007
rect 15151 7973 15160 8007
rect 15108 7964 15160 7973
rect 5540 7828 5592 7880
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 6092 7828 6144 7880
rect 6276 7828 6328 7880
rect 6920 7760 6972 7812
rect 7196 7828 7248 7880
rect 9772 7896 9824 7948
rect 10876 7896 10928 7948
rect 12072 7896 12124 7948
rect 8024 7871 8076 7880
rect 8024 7837 8069 7871
rect 8069 7837 8076 7871
rect 8024 7828 8076 7837
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8392 7871 8444 7880
rect 8392 7837 8402 7871
rect 8402 7837 8436 7871
rect 8436 7837 8444 7871
rect 8392 7828 8444 7837
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9404 7828 9456 7880
rect 9680 7828 9732 7880
rect 10048 7871 10100 7880
rect 10048 7837 10058 7871
rect 10058 7837 10100 7871
rect 10048 7828 10100 7837
rect 10140 7828 10192 7880
rect 10968 7828 11020 7880
rect 7380 7760 7432 7812
rect 7840 7803 7892 7812
rect 7840 7769 7849 7803
rect 7849 7769 7883 7803
rect 7883 7769 7892 7803
rect 7840 7760 7892 7769
rect 4620 7692 4672 7744
rect 4896 7692 4948 7744
rect 9036 7735 9088 7744
rect 9036 7701 9045 7735
rect 9045 7701 9079 7735
rect 9079 7701 9088 7735
rect 9036 7692 9088 7701
rect 10508 7692 10560 7744
rect 10600 7692 10652 7744
rect 12256 7760 12308 7812
rect 14372 7896 14424 7948
rect 16580 7964 16632 8016
rect 17408 7964 17460 8016
rect 17500 8007 17552 8016
rect 17500 7973 17509 8007
rect 17509 7973 17543 8007
rect 17543 7973 17552 8007
rect 17500 7964 17552 7973
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 14832 7828 14884 7880
rect 15568 7871 15620 7880
rect 14556 7760 14608 7812
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 17224 7896 17276 7948
rect 17868 7896 17920 7948
rect 16028 7871 16080 7880
rect 16028 7837 16037 7871
rect 16037 7837 16071 7871
rect 16071 7837 16080 7871
rect 16028 7828 16080 7837
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 16304 7828 16356 7880
rect 15476 7803 15528 7812
rect 15476 7769 15485 7803
rect 15485 7769 15519 7803
rect 15519 7769 15528 7803
rect 15476 7760 15528 7769
rect 16580 7828 16632 7880
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 17500 7828 17552 7880
rect 18420 7871 18472 7880
rect 18420 7837 18429 7871
rect 18429 7837 18463 7871
rect 18463 7837 18472 7871
rect 18420 7828 18472 7837
rect 12348 7692 12400 7744
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 13452 7692 13504 7744
rect 13728 7692 13780 7744
rect 14924 7692 14976 7744
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 16304 7692 16356 7744
rect 16764 7692 16816 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 3332 7488 3384 7540
rect 5816 7488 5868 7540
rect 6736 7488 6788 7540
rect 9036 7488 9088 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 10876 7531 10928 7540
rect 10876 7497 10885 7531
rect 10885 7497 10919 7531
rect 10919 7497 10928 7531
rect 10876 7488 10928 7497
rect 10968 7488 11020 7540
rect 12256 7488 12308 7540
rect 13452 7531 13504 7540
rect 13452 7497 13461 7531
rect 13461 7497 13495 7531
rect 13495 7497 13504 7531
rect 13452 7488 13504 7497
rect 14004 7488 14056 7540
rect 15108 7488 15160 7540
rect 4252 7420 4304 7472
rect 5540 7420 5592 7472
rect 6828 7420 6880 7472
rect 2504 7352 2556 7404
rect 2688 7352 2740 7404
rect 4804 7352 4856 7404
rect 2596 7216 2648 7268
rect 4712 7148 4764 7200
rect 5724 7216 5776 7268
rect 6920 7395 6972 7404
rect 6920 7361 6928 7395
rect 6928 7361 6962 7395
rect 6962 7361 6972 7395
rect 6920 7352 6972 7361
rect 9588 7463 9640 7472
rect 9588 7429 9597 7463
rect 9597 7429 9631 7463
rect 9631 7429 9640 7463
rect 9588 7420 9640 7429
rect 12072 7420 12124 7472
rect 12164 7420 12216 7472
rect 13268 7420 13320 7472
rect 7104 7395 7156 7404
rect 7104 7361 7113 7395
rect 7113 7361 7147 7395
rect 7147 7361 7156 7395
rect 7104 7352 7156 7361
rect 9404 7352 9456 7404
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 7656 7284 7708 7336
rect 12348 7284 12400 7336
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14464 7420 14516 7472
rect 14372 7395 14424 7404
rect 14372 7361 14381 7395
rect 14381 7361 14415 7395
rect 14415 7361 14424 7395
rect 14372 7352 14424 7361
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 14832 7395 14884 7404
rect 14832 7361 14841 7395
rect 14841 7361 14875 7395
rect 14875 7361 14884 7395
rect 14832 7352 14884 7361
rect 14924 7395 14976 7404
rect 14924 7361 14933 7395
rect 14933 7361 14967 7395
rect 14967 7361 14976 7395
rect 14924 7352 14976 7361
rect 17960 7488 18012 7540
rect 17500 7463 17552 7472
rect 17500 7429 17509 7463
rect 17509 7429 17543 7463
rect 17543 7429 17552 7463
rect 17500 7420 17552 7429
rect 17592 7420 17644 7472
rect 7840 7216 7892 7268
rect 11980 7216 12032 7268
rect 13820 7216 13872 7268
rect 14096 7216 14148 7268
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 16764 7395 16816 7404
rect 16764 7361 16773 7395
rect 16773 7361 16807 7395
rect 16807 7361 16816 7395
rect 16764 7352 16816 7361
rect 17132 7352 17184 7404
rect 18052 7284 18104 7336
rect 15476 7216 15528 7268
rect 16120 7216 16172 7268
rect 17132 7216 17184 7268
rect 17224 7216 17276 7268
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 12164 7148 12216 7200
rect 12624 7148 12676 7200
rect 15016 7148 15068 7200
rect 15108 7191 15160 7200
rect 15108 7157 15117 7191
rect 15117 7157 15151 7191
rect 15151 7157 15160 7191
rect 15108 7148 15160 7157
rect 15384 7148 15436 7200
rect 17316 7191 17368 7200
rect 17316 7157 17325 7191
rect 17325 7157 17359 7191
rect 17359 7157 17368 7191
rect 17316 7148 17368 7157
rect 17960 7216 18012 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 5448 6944 5500 6996
rect 6184 6944 6236 6996
rect 11612 6944 11664 6996
rect 9864 6876 9916 6928
rect 12164 6944 12216 6996
rect 12716 6944 12768 6996
rect 4436 6808 4488 6860
rect 7104 6851 7156 6860
rect 7104 6817 7113 6851
rect 7113 6817 7147 6851
rect 7147 6817 7156 6851
rect 7104 6808 7156 6817
rect 6920 6740 6972 6792
rect 8576 6808 8628 6860
rect 8208 6740 8260 6792
rect 10048 6808 10100 6860
rect 16764 6876 16816 6928
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 4528 6715 4580 6724
rect 4528 6681 4537 6715
rect 4537 6681 4571 6715
rect 4571 6681 4580 6715
rect 4528 6672 4580 6681
rect 4804 6672 4856 6724
rect 9588 6672 9640 6724
rect 11612 6851 11664 6860
rect 11612 6817 11621 6851
rect 11621 6817 11655 6851
rect 11655 6817 11664 6851
rect 11612 6808 11664 6817
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 10784 6740 10836 6792
rect 16580 6808 16632 6860
rect 4620 6604 4672 6656
rect 12072 6672 12124 6724
rect 9772 6604 9824 6656
rect 10416 6604 10468 6656
rect 11152 6604 11204 6656
rect 11796 6604 11848 6656
rect 12348 6604 12400 6656
rect 12624 6604 12676 6656
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 17592 6944 17644 6996
rect 17224 6783 17276 6792
rect 17224 6749 17233 6783
rect 17233 6749 17267 6783
rect 17267 6749 17276 6783
rect 17224 6740 17276 6749
rect 17316 6740 17368 6792
rect 18420 6740 18472 6792
rect 13452 6604 13504 6656
rect 15016 6604 15068 6656
rect 16212 6604 16264 6656
rect 17316 6647 17368 6656
rect 17316 6613 17325 6647
rect 17325 6613 17359 6647
rect 17359 6613 17368 6647
rect 17316 6604 17368 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 4528 6400 4580 6452
rect 4436 6307 4488 6316
rect 4436 6273 4445 6307
rect 4445 6273 4479 6307
rect 4479 6273 4488 6307
rect 4436 6264 4488 6273
rect 6920 6400 6972 6452
rect 8116 6400 8168 6452
rect 8760 6400 8812 6452
rect 4804 6196 4856 6248
rect 2964 6060 3016 6112
rect 7932 6332 7984 6384
rect 9312 6400 9364 6452
rect 10784 6400 10836 6452
rect 11612 6400 11664 6452
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7656 6264 7708 6316
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 9956 6332 10008 6384
rect 8852 6307 8904 6316
rect 8852 6273 8861 6307
rect 8861 6273 8895 6307
rect 8895 6273 8904 6307
rect 8852 6264 8904 6273
rect 8944 6264 8996 6316
rect 9772 6264 9824 6316
rect 10048 6307 10100 6316
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10232 6264 10284 6316
rect 10692 6307 10744 6316
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 11980 6332 12032 6384
rect 13820 6400 13872 6452
rect 15936 6400 15988 6452
rect 13452 6332 13504 6384
rect 15476 6332 15528 6384
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 11520 6307 11572 6316
rect 11520 6273 11529 6307
rect 11529 6273 11563 6307
rect 11563 6273 11572 6307
rect 11520 6264 11572 6273
rect 14832 6264 14884 6316
rect 10784 6196 10836 6248
rect 10876 6196 10928 6248
rect 12532 6196 12584 6248
rect 14556 6196 14608 6248
rect 15108 6196 15160 6248
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 15568 6196 15620 6248
rect 16212 6307 16264 6316
rect 16212 6273 16221 6307
rect 16221 6273 16255 6307
rect 16255 6273 16264 6307
rect 16212 6264 16264 6273
rect 16304 6307 16356 6316
rect 16304 6273 16313 6307
rect 16313 6273 16347 6307
rect 16347 6273 16356 6307
rect 16304 6264 16356 6273
rect 16488 6307 16540 6316
rect 16488 6273 16497 6307
rect 16497 6273 16531 6307
rect 16531 6273 16540 6307
rect 16488 6264 16540 6273
rect 17408 6307 17460 6316
rect 17408 6273 17417 6307
rect 17417 6273 17451 6307
rect 17451 6273 17460 6307
rect 17408 6264 17460 6273
rect 16396 6196 16448 6248
rect 16580 6196 16632 6248
rect 17224 6196 17276 6248
rect 17500 6196 17552 6248
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 8024 6171 8076 6180
rect 8024 6137 8033 6171
rect 8033 6137 8067 6171
rect 8067 6137 8076 6171
rect 8024 6128 8076 6137
rect 8852 6128 8904 6180
rect 9864 6128 9916 6180
rect 10048 6128 10100 6180
rect 10600 6128 10652 6180
rect 7288 6060 7340 6112
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 8668 6060 8720 6112
rect 8760 6060 8812 6112
rect 10140 6060 10192 6112
rect 10508 6060 10560 6112
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 16028 6128 16080 6180
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 15752 6060 15804 6112
rect 15844 6060 15896 6112
rect 16764 6060 16816 6112
rect 17316 6060 17368 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 5264 5856 5316 5908
rect 9128 5856 9180 5908
rect 4804 5788 4856 5840
rect 5356 5788 5408 5840
rect 7472 5788 7524 5840
rect 7748 5788 7800 5840
rect 9036 5788 9088 5840
rect 7288 5695 7340 5704
rect 7288 5661 7297 5695
rect 7297 5661 7331 5695
rect 7331 5661 7340 5695
rect 7288 5652 7340 5661
rect 7748 5652 7800 5704
rect 8852 5720 8904 5772
rect 4896 5584 4948 5636
rect 8208 5652 8260 5704
rect 9864 5856 9916 5908
rect 10140 5788 10192 5840
rect 10968 5856 11020 5908
rect 11980 5899 12032 5908
rect 11980 5865 11989 5899
rect 11989 5865 12023 5899
rect 12023 5865 12032 5899
rect 11980 5856 12032 5865
rect 15200 5856 15252 5908
rect 15568 5856 15620 5908
rect 16212 5856 16264 5908
rect 9312 5695 9364 5704
rect 9312 5661 9321 5695
rect 9321 5661 9355 5695
rect 9355 5661 9364 5695
rect 9312 5652 9364 5661
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 8300 5584 8352 5636
rect 8392 5627 8444 5636
rect 8392 5593 8401 5627
rect 8401 5593 8435 5627
rect 8435 5593 8444 5627
rect 8392 5584 8444 5593
rect 8760 5584 8812 5636
rect 9956 5652 10008 5704
rect 10324 5652 10376 5704
rect 9680 5584 9732 5636
rect 10048 5584 10100 5636
rect 10876 5720 10928 5772
rect 12348 5720 12400 5772
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 12072 5652 12124 5704
rect 12716 5695 12768 5704
rect 12716 5661 12725 5695
rect 12725 5661 12759 5695
rect 12759 5661 12768 5695
rect 12716 5652 12768 5661
rect 12256 5584 12308 5636
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 15200 5763 15252 5772
rect 15200 5729 15209 5763
rect 15209 5729 15243 5763
rect 15243 5729 15252 5763
rect 15200 5720 15252 5729
rect 16396 5788 16448 5840
rect 15660 5720 15712 5772
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 15384 5652 15436 5704
rect 15936 5652 15988 5704
rect 16120 5695 16172 5704
rect 16120 5661 16132 5695
rect 16132 5661 16166 5695
rect 16166 5661 16172 5695
rect 17040 5856 17092 5908
rect 16120 5652 16172 5661
rect 16580 5695 16632 5704
rect 16580 5661 16589 5695
rect 16589 5661 16623 5695
rect 16623 5661 16632 5695
rect 16580 5652 16632 5661
rect 16764 5695 16816 5704
rect 16764 5661 16773 5695
rect 16773 5661 16807 5695
rect 16807 5661 16816 5695
rect 16764 5652 16816 5661
rect 17316 5652 17368 5704
rect 18604 5652 18656 5704
rect 8116 5516 8168 5568
rect 8484 5516 8536 5568
rect 8668 5516 8720 5568
rect 9128 5516 9180 5568
rect 10784 5516 10836 5568
rect 10876 5559 10928 5568
rect 10876 5525 10885 5559
rect 10885 5525 10919 5559
rect 10919 5525 10928 5559
rect 10876 5516 10928 5525
rect 12164 5516 12216 5568
rect 14648 5584 14700 5636
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 16856 5627 16908 5636
rect 16856 5593 16865 5627
rect 16865 5593 16899 5627
rect 16899 5593 16908 5627
rect 16856 5584 16908 5593
rect 17132 5559 17184 5568
rect 17132 5525 17141 5559
rect 17141 5525 17175 5559
rect 17175 5525 17184 5559
rect 17132 5516 17184 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 10232 5312 10284 5364
rect 5356 5176 5408 5228
rect 5540 5244 5592 5296
rect 8300 5244 8352 5296
rect 9496 5244 9548 5296
rect 9956 5287 10008 5296
rect 9956 5253 9965 5287
rect 9965 5253 9999 5287
rect 9999 5253 10008 5287
rect 9956 5244 10008 5253
rect 7932 5176 7984 5228
rect 8484 5176 8536 5228
rect 8760 5176 8812 5228
rect 8944 5219 8996 5228
rect 8944 5185 8953 5219
rect 8953 5185 8987 5219
rect 8987 5185 8996 5219
rect 8944 5176 8996 5185
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 9404 5176 9456 5228
rect 8392 5108 8444 5160
rect 9588 5108 9640 5160
rect 9036 5040 9088 5092
rect 10140 5176 10192 5228
rect 10876 5312 10928 5364
rect 15752 5312 15804 5364
rect 16120 5312 16172 5364
rect 16488 5312 16540 5364
rect 12164 5244 12216 5296
rect 13636 5244 13688 5296
rect 14648 5287 14700 5296
rect 14648 5253 14657 5287
rect 14657 5253 14691 5287
rect 14691 5253 14700 5287
rect 14648 5244 14700 5253
rect 10692 5176 10744 5228
rect 12256 5176 12308 5228
rect 12532 5176 12584 5228
rect 14832 5219 14884 5228
rect 14832 5185 14841 5219
rect 14841 5185 14875 5219
rect 14875 5185 14884 5219
rect 14832 5176 14884 5185
rect 15476 5244 15528 5296
rect 15200 5219 15252 5228
rect 15200 5185 15209 5219
rect 15209 5185 15243 5219
rect 15243 5185 15252 5219
rect 15200 5176 15252 5185
rect 16856 5244 16908 5296
rect 16028 5176 16080 5228
rect 17132 5176 17184 5228
rect 16212 5108 16264 5160
rect 4712 4972 4764 5024
rect 5264 4972 5316 5024
rect 16304 5040 16356 5092
rect 14464 4972 14516 5024
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 5540 4768 5592 4820
rect 5908 4811 5960 4820
rect 5908 4777 5917 4811
rect 5917 4777 5951 4811
rect 5951 4777 5960 4811
rect 5908 4768 5960 4777
rect 6644 4768 6696 4820
rect 9036 4811 9088 4820
rect 9036 4777 9045 4811
rect 9045 4777 9079 4811
rect 9079 4777 9088 4811
rect 9036 4768 9088 4777
rect 9312 4768 9364 4820
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 4528 4632 4580 4684
rect 9404 4700 9456 4752
rect 5540 4564 5592 4616
rect 5816 4564 5868 4616
rect 6828 4564 6880 4616
rect 8760 4564 8812 4616
rect 9128 4632 9180 4684
rect 9036 4564 9088 4616
rect 12348 4564 12400 4616
rect 12624 4564 12676 4616
rect 4436 4539 4488 4548
rect 4436 4505 4445 4539
rect 4445 4505 4479 4539
rect 4479 4505 4488 4539
rect 4436 4496 4488 4505
rect 6644 4539 6696 4548
rect 6644 4505 6653 4539
rect 6653 4505 6687 4539
rect 6687 4505 6696 4539
rect 6644 4496 6696 4505
rect 6368 4471 6420 4480
rect 6368 4437 6377 4471
rect 6377 4437 6411 4471
rect 6411 4437 6420 4471
rect 6368 4428 6420 4437
rect 6460 4428 6512 4480
rect 12348 4471 12400 4480
rect 12348 4437 12357 4471
rect 12357 4437 12391 4471
rect 12391 4437 12400 4471
rect 12348 4428 12400 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4436 4224 4488 4276
rect 4620 4224 4672 4276
rect 4712 4199 4764 4208
rect 4712 4165 4721 4199
rect 4721 4165 4755 4199
rect 4755 4165 4764 4199
rect 4712 4156 4764 4165
rect 5816 4199 5868 4208
rect 5816 4165 5825 4199
rect 5825 4165 5859 4199
rect 5859 4165 5868 4199
rect 5816 4156 5868 4165
rect 5264 4088 5316 4140
rect 5448 4088 5500 4140
rect 8760 4224 8812 4276
rect 9404 4224 9456 4276
rect 12256 4224 12308 4276
rect 6460 4088 6512 4140
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 10508 4199 10560 4208
rect 10508 4165 10517 4199
rect 10517 4165 10551 4199
rect 10551 4165 10560 4199
rect 10508 4156 10560 4165
rect 11060 4156 11112 4208
rect 13820 4156 13872 4208
rect 9220 4088 9272 4140
rect 9680 4088 9732 4140
rect 9956 4088 10008 4140
rect 10692 4088 10744 4140
rect 11704 4088 11756 4140
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 12164 4131 12216 4140
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 8208 4020 8260 4072
rect 12164 4097 12173 4131
rect 12173 4097 12207 4131
rect 12207 4097 12216 4131
rect 12164 4088 12216 4097
rect 12348 4131 12400 4140
rect 12348 4097 12357 4131
rect 12357 4097 12391 4131
rect 12391 4097 12400 4131
rect 12348 4088 12400 4097
rect 12072 4020 12124 4072
rect 10140 3995 10192 4004
rect 10140 3961 10149 3995
rect 10149 3961 10183 3995
rect 10183 3961 10192 3995
rect 10140 3952 10192 3961
rect 10416 3952 10468 4004
rect 12624 4088 12676 4140
rect 12624 3952 12676 4004
rect 4804 3884 4856 3936
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 5908 3884 5960 3936
rect 6184 3927 6236 3936
rect 6184 3893 6193 3927
rect 6193 3893 6227 3927
rect 6227 3893 6236 3927
rect 6184 3884 6236 3893
rect 10600 3884 10652 3936
rect 14556 3884 14608 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 5540 3680 5592 3732
rect 4804 3612 4856 3664
rect 6184 3655 6236 3664
rect 6184 3621 6193 3655
rect 6193 3621 6227 3655
rect 6227 3621 6236 3655
rect 6184 3612 6236 3621
rect 6828 3680 6880 3732
rect 7012 3612 7064 3664
rect 8208 3612 8260 3664
rect 9404 3612 9456 3664
rect 10140 3680 10192 3732
rect 11888 3680 11940 3732
rect 12348 3680 12400 3732
rect 6368 3544 6420 3596
rect 8852 3476 8904 3528
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 11704 3544 11756 3596
rect 5724 3408 5776 3460
rect 6920 3408 6972 3460
rect 8116 3408 8168 3460
rect 8208 3408 8260 3460
rect 9680 3451 9732 3460
rect 9680 3417 9689 3451
rect 9689 3417 9723 3451
rect 9723 3417 9732 3451
rect 9680 3408 9732 3417
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 11520 3476 11572 3528
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 13636 3476 13688 3528
rect 13820 3723 13872 3732
rect 13820 3689 13829 3723
rect 13829 3689 13863 3723
rect 13863 3689 13872 3723
rect 13820 3680 13872 3689
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 8852 3340 8904 3392
rect 14832 3408 14884 3460
rect 11060 3340 11112 3392
rect 12072 3340 12124 3392
rect 13544 3383 13596 3392
rect 13544 3349 13553 3383
rect 13553 3349 13587 3383
rect 13587 3349 13596 3383
rect 13544 3340 13596 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 8024 3068 8076 3120
rect 6552 3000 6604 3052
rect 10140 3136 10192 3188
rect 12532 3136 12584 3188
rect 14832 3136 14884 3188
rect 8852 3111 8904 3120
rect 8852 3077 8861 3111
rect 8861 3077 8895 3111
rect 8895 3077 8904 3111
rect 8852 3068 8904 3077
rect 10416 3068 10468 3120
rect 10508 3111 10560 3120
rect 10508 3077 10517 3111
rect 10517 3077 10551 3111
rect 10551 3077 10560 3111
rect 10508 3068 10560 3077
rect 7104 2932 7156 2984
rect 8944 2932 8996 2984
rect 9220 2932 9272 2984
rect 10692 3043 10744 3052
rect 10692 3009 10701 3043
rect 10701 3009 10735 3043
rect 10735 3009 10744 3043
rect 10692 3000 10744 3009
rect 11060 3000 11112 3052
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11520 3068 11572 3120
rect 12348 3068 12400 3120
rect 12072 3043 12124 3052
rect 12072 3009 12081 3043
rect 12081 3009 12115 3043
rect 12115 3009 12124 3043
rect 12072 3000 12124 3009
rect 14004 3068 14056 3120
rect 8116 2796 8168 2848
rect 9220 2796 9272 2848
rect 9404 2796 9456 2848
rect 10600 2796 10652 2848
rect 13544 2796 13596 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 7104 2592 7156 2644
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 8668 2635 8720 2644
rect 8668 2601 8677 2635
rect 8677 2601 8711 2635
rect 8711 2601 8720 2635
rect 8668 2592 8720 2601
rect 14004 2592 14056 2644
rect 6368 2524 6420 2576
rect 8484 2524 8536 2576
rect 9772 2524 9824 2576
rect 8116 2431 8168 2440
rect 8116 2397 8125 2431
rect 8125 2397 8159 2431
rect 8159 2397 8168 2431
rect 8116 2388 8168 2397
rect 7196 2320 7248 2372
rect 7748 2320 7800 2372
rect 8392 2388 8444 2440
rect 9680 2388 9732 2440
rect 13636 2431 13688 2440
rect 13636 2397 13645 2431
rect 13645 2397 13679 2431
rect 13679 2397 13688 2431
rect 13636 2388 13688 2397
rect 9036 2320 9088 2372
rect 8760 2252 8812 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5814 21382 5870 22182
rect 6458 21382 6514 22182
rect 12898 21382 12954 22182
rect 13542 21382 13598 22182
rect 13648 21406 13860 21434
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5828 19310 5856 21382
rect 6472 19378 6500 21382
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6184 19372 6236 19378
rect 6184 19314 6236 19320
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 5816 19304 5868 19310
rect 5816 19246 5868 19252
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4620 18760 4672 18766
rect 4672 18708 4752 18714
rect 4620 18702 4752 18708
rect 4344 18692 4396 18698
rect 4632 18686 4752 18702
rect 4344 18634 4396 18640
rect 4356 18290 4384 18634
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4632 18358 4660 18566
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4344 18284 4396 18290
rect 4344 18226 4396 18232
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 1412 17785 1440 18158
rect 4724 18086 4752 18686
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2504 17536 2556 17542
rect 2504 17478 2556 17484
rect 2424 17338 2452 17478
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 1768 17264 1820 17270
rect 1768 17206 1820 17212
rect 1676 16516 1728 16522
rect 1676 16458 1728 16464
rect 848 16108 900 16114
rect 848 16050 900 16056
rect 860 15881 888 16050
rect 846 15872 902 15881
rect 846 15807 902 15816
rect 1688 15502 1716 16458
rect 1780 16250 1808 17206
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1964 16590 1992 16934
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1860 16448 1912 16454
rect 1860 16390 1912 16396
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1780 15570 1808 16186
rect 1872 16114 1900 16390
rect 2332 16250 2360 17138
rect 2424 16998 2452 17274
rect 2516 17270 2544 17478
rect 2504 17264 2556 17270
rect 2504 17206 2556 17212
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2608 16794 2636 17818
rect 4068 17808 4120 17814
rect 4068 17750 4120 17756
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2596 16788 2648 16794
rect 2648 16748 2728 16776
rect 2596 16730 2648 16736
rect 2596 16448 2648 16454
rect 2596 16390 2648 16396
rect 2320 16244 2372 16250
rect 2320 16186 2372 16192
rect 1860 16108 1912 16114
rect 1860 16050 1912 16056
rect 2608 16046 2636 16390
rect 2700 16182 2728 16748
rect 2792 16522 2820 17614
rect 2884 16590 2912 17682
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 3160 17338 3188 17614
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 3056 17196 3108 17202
rect 2976 17156 3056 17184
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2688 16176 2740 16182
rect 2688 16118 2740 16124
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 1768 15564 1820 15570
rect 1768 15506 1820 15512
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1688 15162 1716 15438
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 848 15020 900 15026
rect 848 14962 900 14968
rect 860 14929 888 14962
rect 1780 14958 1808 15506
rect 1676 14952 1728 14958
rect 846 14920 902 14929
rect 1676 14894 1728 14900
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 846 14855 902 14864
rect 1688 14550 1716 14894
rect 2228 14884 2280 14890
rect 2228 14826 2280 14832
rect 2240 14618 2268 14826
rect 2228 14612 2280 14618
rect 2228 14554 2280 14560
rect 1676 14544 1728 14550
rect 846 14512 902 14521
rect 1676 14486 1728 14492
rect 2044 14544 2096 14550
rect 2044 14486 2096 14492
rect 846 14447 902 14456
rect 860 14414 888 14447
rect 848 14408 900 14414
rect 848 14350 900 14356
rect 2056 13938 2084 14486
rect 2240 14482 2268 14554
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2608 13938 2636 15982
rect 2700 15502 2728 16118
rect 2872 15564 2924 15570
rect 2872 15506 2924 15512
rect 2688 15496 2740 15502
rect 2688 15438 2740 15444
rect 2884 15026 2912 15506
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2976 14618 3004 17156
rect 3056 17138 3108 17144
rect 3160 16794 3188 17274
rect 3988 17270 4016 17682
rect 4080 17338 4108 17750
rect 4068 17332 4120 17338
rect 4068 17274 4120 17280
rect 3976 17264 4028 17270
rect 3976 17206 4028 17212
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3148 16788 3200 16794
rect 3148 16730 3200 16736
rect 3252 15910 3280 17138
rect 4620 17128 4672 17134
rect 4620 17070 4672 17076
rect 3332 16992 3384 16998
rect 3332 16934 3384 16940
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3344 15026 3372 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16590 4660 17070
rect 4724 16998 4752 18022
rect 5276 17882 5304 18634
rect 5644 18426 5672 19178
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5724 18828 5776 18834
rect 5724 18770 5776 18776
rect 5632 18420 5684 18426
rect 5632 18362 5684 18368
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5368 18086 5396 18158
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 5368 17746 5396 18022
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 5368 17338 5396 17682
rect 5736 17542 5764 18770
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4712 16992 4764 16998
rect 4712 16934 4764 16940
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3712 15026 3740 15846
rect 3896 15026 3924 15914
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4160 15632 4212 15638
rect 4160 15574 4212 15580
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3516 15020 3568 15026
rect 3516 14962 3568 14968
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3056 14816 3108 14822
rect 3056 14758 3108 14764
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3068 14482 3096 14758
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2056 13394 2084 13874
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 2148 13326 2176 13874
rect 2596 13728 2648 13734
rect 2596 13670 2648 13676
rect 2608 13462 2636 13670
rect 2596 13456 2648 13462
rect 2596 13398 2648 13404
rect 3332 13456 3384 13462
rect 3332 13398 3384 13404
rect 2688 13388 2740 13394
rect 2688 13330 2740 13336
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 848 13184 900 13190
rect 846 13152 848 13161
rect 900 13152 902 13161
rect 846 13087 902 13096
rect 848 12232 900 12238
rect 846 12200 848 12209
rect 900 12200 902 12209
rect 846 12135 902 12144
rect 846 11792 902 11801
rect 846 11727 848 11736
rect 900 11727 902 11736
rect 848 11698 900 11704
rect 1412 11354 1440 13262
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 1584 12708 1636 12714
rect 1584 12650 1636 12656
rect 1596 12442 1624 12650
rect 1676 12640 1728 12646
rect 1676 12582 1728 12588
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1688 12306 1716 12582
rect 1676 12300 1728 12306
rect 1676 12242 1728 12248
rect 2056 11898 2084 12786
rect 2148 12646 2176 13262
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12782 2268 13126
rect 2700 12782 2728 13330
rect 3344 13326 3372 13398
rect 3528 13326 3556 14962
rect 3608 14952 3660 14958
rect 3608 14894 3660 14900
rect 3620 14346 3648 14894
rect 3896 14618 3924 14962
rect 4172 14906 4200 15574
rect 4356 15502 4384 15642
rect 4632 15570 4660 16390
rect 4724 16028 4752 16934
rect 4816 16182 4844 17138
rect 5368 16726 5396 17274
rect 5736 17202 5764 17478
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5540 16788 5592 16794
rect 5736 16776 5764 17138
rect 5592 16748 5764 16776
rect 5540 16730 5592 16736
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5368 16590 5396 16662
rect 5736 16590 5764 16748
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5724 16584 5776 16590
rect 5724 16526 5776 16532
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5368 16182 5396 16390
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 5356 16176 5408 16182
rect 5356 16118 5408 16124
rect 5736 16114 5764 16526
rect 5724 16108 5776 16114
rect 5724 16050 5776 16056
rect 4896 16040 4948 16046
rect 4724 16000 4896 16028
rect 4896 15982 4948 15988
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4620 15564 4672 15570
rect 4620 15506 4672 15512
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4356 15162 4384 15438
rect 4528 15428 4580 15434
rect 4528 15370 4580 15376
rect 4344 15156 4396 15162
rect 4344 15098 4396 15104
rect 4540 15026 4568 15370
rect 4632 15094 4660 15506
rect 4816 15502 4844 15846
rect 4908 15638 4936 15982
rect 4896 15632 4948 15638
rect 4896 15574 4948 15580
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 3988 14878 4200 14906
rect 4252 14952 4304 14958
rect 4304 14912 4476 14940
rect 4252 14894 4304 14900
rect 4448 14906 4476 14912
rect 4448 14890 4568 14906
rect 4448 14884 4580 14890
rect 4448 14878 4528 14884
rect 3988 14618 4016 14878
rect 4528 14826 4580 14832
rect 4724 14822 4752 15438
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3608 14340 3660 14346
rect 3608 14282 3660 14288
rect 3896 13326 3924 14350
rect 3976 14272 4028 14278
rect 3976 14214 4028 14220
rect 3988 13394 4016 14214
rect 3976 13388 4028 13394
rect 3976 13330 4028 13336
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2688 12776 2740 12782
rect 2688 12718 2740 12724
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2240 12238 2268 12718
rect 2872 12640 2924 12646
rect 2700 12600 2872 12628
rect 2700 12434 2728 12600
rect 2872 12582 2924 12588
rect 2608 12406 2728 12434
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2516 12170 2544 12310
rect 2608 12238 2636 12406
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2044 11892 2096 11898
rect 2044 11834 2096 11840
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1596 10810 1624 11630
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 11082 2176 11494
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 860 10441 888 10610
rect 846 10432 902 10441
rect 846 10367 902 10376
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1596 9450 1624 10746
rect 2608 10606 2636 12174
rect 2976 12102 3004 12718
rect 3068 12714 3096 13262
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3252 12986 3280 13194
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 3056 12708 3108 12714
rect 3056 12650 3108 12656
rect 3804 12442 3832 12786
rect 3896 12782 3924 13262
rect 3976 13184 4028 13190
rect 3976 13126 4028 13132
rect 3988 12850 4016 13126
rect 4080 12850 4108 14758
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4632 14618 4660 14758
rect 4816 14618 4844 15438
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4908 14498 4936 14894
rect 5092 14618 5120 14894
rect 5264 14884 5316 14890
rect 5264 14826 5316 14832
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4816 14470 4936 14498
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4160 13252 4212 13258
rect 4160 13194 4212 13200
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3884 12776 3936 12782
rect 4172 12730 4200 13194
rect 4632 12986 4660 14418
rect 4816 14414 4844 14470
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4816 13530 4844 14350
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 3884 12718 3936 12724
rect 4080 12714 4200 12730
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 3976 12708 4028 12714
rect 3976 12650 4028 12656
rect 4068 12708 4200 12714
rect 4120 12702 4200 12708
rect 4068 12650 4120 12656
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3424 12368 3476 12374
rect 3424 12310 3476 12316
rect 3436 12238 3464 12310
rect 3988 12238 4016 12650
rect 4080 12288 4108 12650
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4160 12300 4212 12306
rect 4080 12260 4160 12288
rect 4160 12242 4212 12248
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2700 10674 2728 11834
rect 3436 11150 3464 12174
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11150 4016 12038
rect 4448 11898 4476 12174
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4632 11778 4660 12718
rect 4724 12238 4752 12786
rect 4988 12776 5040 12782
rect 4988 12718 5040 12724
rect 5000 12238 5028 12718
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4988 12232 5040 12238
rect 4988 12174 5040 12180
rect 5276 12102 5304 14826
rect 5368 12442 5396 15302
rect 5828 15094 5856 18906
rect 6104 18358 6132 19314
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 6196 18290 6224 19314
rect 6644 19304 6696 19310
rect 6644 19246 6696 19252
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6472 18426 6500 18702
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6184 18284 6236 18290
rect 6184 18226 6236 18232
rect 6184 17876 6236 17882
rect 6184 17818 6236 17824
rect 6196 17338 6224 17818
rect 6276 17672 6328 17678
rect 6276 17614 6328 17620
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6092 17196 6144 17202
rect 6092 17138 6144 17144
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6012 16454 6040 16526
rect 6104 16454 6132 17138
rect 6288 16794 6316 17614
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6288 16590 6316 16730
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6276 16448 6328 16454
rect 6276 16390 6328 16396
rect 6012 15978 6040 16390
rect 6104 16250 6132 16390
rect 6092 16244 6144 16250
rect 6092 16186 6144 16192
rect 6288 16114 6316 16390
rect 6472 16182 6500 17478
rect 6656 16658 6684 19246
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 6748 17202 6776 18566
rect 7024 17270 7052 19382
rect 11336 19372 11388 19378
rect 11336 19314 11388 19320
rect 9312 19236 9364 19242
rect 9312 19178 9364 19184
rect 8022 18320 8078 18329
rect 7748 18284 7800 18290
rect 8022 18255 8078 18264
rect 7748 18226 7800 18232
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7116 17270 7144 17478
rect 7760 17338 7788 18226
rect 7748 17332 7800 17338
rect 7748 17274 7800 17280
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6460 16176 6512 16182
rect 6460 16118 6512 16124
rect 6276 16108 6328 16114
rect 6276 16050 6328 16056
rect 6000 15972 6052 15978
rect 6000 15914 6052 15920
rect 6012 15706 6040 15914
rect 6000 15700 6052 15706
rect 6000 15642 6052 15648
rect 6288 15502 6316 16050
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6092 15360 6144 15366
rect 6092 15302 6144 15308
rect 5816 15088 5868 15094
rect 5816 15030 5868 15036
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 5828 14550 5856 15030
rect 6012 14618 6040 15030
rect 6104 14822 6132 15302
rect 6092 14816 6144 14822
rect 6092 14758 6144 14764
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 5816 14544 5868 14550
rect 5816 14486 5868 14492
rect 6288 14414 6316 15438
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6380 14822 6408 15370
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6380 14550 6408 14758
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5460 12322 5488 14282
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 5828 14074 5856 14214
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5724 13932 5776 13938
rect 5724 13874 5776 13880
rect 5736 13258 5764 13874
rect 5828 13530 5856 14010
rect 6288 14006 6316 14350
rect 6380 14074 6408 14486
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6276 14000 6328 14006
rect 6276 13942 6328 13948
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13530 6408 13670
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5644 12986 5672 13194
rect 5736 12986 5764 13194
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5828 12850 5856 13466
rect 6472 13410 6500 16118
rect 6656 15910 6684 16390
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6748 15094 6776 17138
rect 7760 16114 7788 17274
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 7656 15904 7708 15910
rect 7656 15846 7708 15852
rect 6932 15570 6960 15846
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 7668 15434 7696 15846
rect 7656 15428 7708 15434
rect 7656 15370 7708 15376
rect 6736 15088 6788 15094
rect 6736 15030 6788 15036
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 6748 14618 6776 15030
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6748 14006 6776 14554
rect 7668 14074 7696 15030
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6564 13530 6592 13874
rect 6552 13524 6604 13530
rect 6552 13466 6604 13472
rect 6380 13382 6500 13410
rect 6644 13388 6696 13394
rect 6380 13190 6408 13382
rect 6748 13376 6776 13942
rect 7760 13938 7788 16050
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 6696 13348 6776 13376
rect 6644 13330 6696 13336
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 5920 12986 5948 13126
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6380 12918 6408 13126
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 5540 12844 5592 12850
rect 5540 12786 5592 12792
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5368 12306 5488 12322
rect 5356 12300 5488 12306
rect 5408 12294 5488 12300
rect 5356 12242 5408 12248
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4068 11756 4120 11762
rect 4632 11750 4752 11778
rect 4068 11698 4120 11704
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4080 11082 4108 11698
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4632 11150 4660 11630
rect 4252 11144 4304 11150
rect 4252 11086 4304 11092
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4068 11076 4120 11082
rect 4068 11018 4120 11024
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4172 10674 4200 10950
rect 4264 10810 4292 11086
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 2688 10668 2740 10674
rect 2688 10610 2740 10616
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 2596 10600 2648 10606
rect 2596 10542 2648 10548
rect 2608 10130 2636 10542
rect 2700 10266 2728 10610
rect 3884 10600 3936 10606
rect 4264 10554 4292 10746
rect 4448 10588 4476 11086
rect 4724 10742 4752 11750
rect 5368 11354 5396 12242
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11898 5488 12038
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5552 11558 5580 12786
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4712 10736 4764 10742
rect 4712 10678 4764 10684
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4528 10600 4580 10606
rect 4448 10560 4528 10588
rect 3884 10542 3936 10548
rect 2688 10260 2740 10266
rect 2688 10202 2740 10208
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9586 1716 9862
rect 1872 9586 1900 10066
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 1964 9722 1992 9998
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1964 9586 1992 9658
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1952 9580 2004 9586
rect 1952 9522 2004 9528
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 846 9072 902 9081
rect 846 9007 902 9016
rect 860 8974 888 9007
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 1872 8498 1900 9522
rect 2228 9444 2280 9450
rect 2228 9386 2280 9392
rect 2240 9042 2268 9386
rect 2320 9376 2372 9382
rect 2320 9318 2372 9324
rect 2332 9042 2360 9318
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 2320 9036 2372 9042
rect 2320 8978 2372 8984
rect 2136 8968 2188 8974
rect 2134 8936 2136 8945
rect 2188 8936 2190 8945
rect 2134 8871 2190 8880
rect 2332 8634 2360 8978
rect 2792 8974 2820 9998
rect 3896 9518 3924 10542
rect 4080 10526 4292 10554
rect 4528 10542 4580 10548
rect 4080 10248 4108 10526
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4080 10220 4200 10248
rect 4172 9602 4200 10220
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4080 9586 4200 9602
rect 4068 9580 4200 9586
rect 4120 9574 4200 9580
rect 4068 9522 4120 9528
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 3884 9512 3936 9518
rect 3884 9454 3936 9460
rect 2976 9110 3004 9454
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 1412 8265 1440 8366
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 2516 7886 2544 8434
rect 2608 7954 2636 8774
rect 2792 8430 2820 8910
rect 3160 8906 3188 9318
rect 3896 9178 3924 9454
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3068 8566 3096 8842
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 3240 8356 3292 8362
rect 3240 8298 3292 8304
rect 2688 8288 2740 8294
rect 2688 8230 2740 8236
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2596 7948 2648 7954
rect 2596 7890 2648 7896
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 2516 7410 2544 7822
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2608 7274 2636 7890
rect 2700 7818 2728 8230
rect 2976 7954 3004 8230
rect 2964 7948 3016 7954
rect 2964 7890 3016 7896
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2700 7410 2728 7754
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2976 6118 3004 7890
rect 3252 7886 3280 8298
rect 3344 8294 3372 9114
rect 3516 9036 3568 9042
rect 3568 8996 3648 9024
rect 3516 8978 3568 8984
rect 3620 8566 3648 8996
rect 3988 8974 4016 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9042 4660 9862
rect 4724 9654 4752 9998
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 3792 8968 3844 8974
rect 3792 8910 3844 8916
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 3608 8560 3660 8566
rect 3804 8537 3832 8910
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3608 8502 3660 8508
rect 3790 8528 3846 8537
rect 3790 8463 3792 8472
rect 3844 8463 3846 8472
rect 3792 8434 3844 8440
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3988 7886 4016 8774
rect 4356 8634 4384 8910
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4724 8498 4752 9318
rect 4816 8974 4844 10610
rect 5368 10470 5396 11086
rect 5552 10810 5580 11290
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5448 10736 5500 10742
rect 5448 10678 5500 10684
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4908 8820 4936 8978
rect 5092 8906 5120 9046
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4816 8792 4936 8820
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4172 8276 4200 8434
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4080 8248 4200 8276
rect 4540 8276 4568 8366
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4540 8248 4660 8276
rect 4080 8090 4108 8248
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8090 4660 8248
rect 4068 8084 4120 8090
rect 4068 8026 4120 8032
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4724 7954 4752 8298
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3344 7546 3372 7822
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 4264 7478 4292 7754
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4252 7472 4304 7478
rect 4252 7414 4304 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6984 4660 7686
rect 4816 7410 4844 8792
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 4908 8362 4936 8570
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4908 7886 4936 8298
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 5184 7834 5212 8570
rect 5276 8498 5304 10406
rect 5368 10266 5396 10406
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 5460 9178 5488 10678
rect 5644 9654 5672 11018
rect 5920 10742 5948 12582
rect 6656 12434 6684 13330
rect 7760 12850 7788 13874
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7944 12986 7972 13194
rect 7932 12980 7984 12986
rect 7932 12922 7984 12928
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6472 12406 6684 12434
rect 6472 12238 6500 12406
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6472 11218 6500 12174
rect 6932 12102 6960 12582
rect 7208 12442 7236 12786
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7944 12306 7972 12786
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 7944 11830 7972 12242
rect 8036 11830 8064 18255
rect 9324 17202 9352 19178
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 9864 18964 9916 18970
rect 9864 18906 9916 18912
rect 9876 18290 9904 18906
rect 10784 18828 10836 18834
rect 10784 18770 10836 18776
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10244 18426 10272 18634
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9508 17610 9536 18022
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9048 15162 9076 16118
rect 9140 15434 9168 16458
rect 9128 15428 9180 15434
rect 9128 15370 9180 15376
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 7932 11824 7984 11830
rect 7932 11766 7984 11772
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6552 11212 6604 11218
rect 6552 11154 6604 11160
rect 6564 10742 6592 11154
rect 7944 11150 7972 11766
rect 8588 11286 8616 15098
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8680 14550 8708 14758
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8680 14006 8708 14486
rect 8668 14000 8720 14006
rect 8668 13942 8720 13948
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 8668 13728 8720 13734
rect 8668 13670 8720 13676
rect 8680 13530 8708 13670
rect 8668 13524 8720 13530
rect 8668 13466 8720 13472
rect 9140 12986 9168 13942
rect 9220 13728 9272 13734
rect 9220 13670 9272 13676
rect 9232 13258 9260 13670
rect 9220 13252 9272 13258
rect 9220 13194 9272 13200
rect 9128 12980 9180 12986
rect 9128 12922 9180 12928
rect 9324 12434 9352 17138
rect 9876 16998 9904 18226
rect 10508 17876 10560 17882
rect 10508 17818 10560 17824
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9508 15706 9536 15982
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9600 14346 9628 14962
rect 9784 14822 9812 15370
rect 9876 14958 9904 16934
rect 9968 16454 9996 17138
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 16046 9996 16390
rect 10060 16114 10088 17682
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10336 17270 10364 17478
rect 10520 17338 10548 17818
rect 10704 17626 10732 18226
rect 10796 17746 10824 18770
rect 11256 18698 11284 19110
rect 11348 18970 11376 19314
rect 12912 19310 12940 21382
rect 13556 21298 13584 21382
rect 13648 21298 13676 21406
rect 13556 21270 13676 21298
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 11336 18964 11388 18970
rect 11336 18906 11388 18912
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11520 18352 11572 18358
rect 11520 18294 11572 18300
rect 11152 18284 11204 18290
rect 11152 18226 11204 18232
rect 11164 18034 11192 18226
rect 11244 18080 11296 18086
rect 11164 18028 11244 18034
rect 11164 18022 11296 18028
rect 11164 18006 11284 18022
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10612 17610 10732 17626
rect 11164 17610 11192 18006
rect 11532 17678 11560 18294
rect 11716 18222 11744 18566
rect 12084 18426 12112 18634
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13096 18426 13124 18566
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 11888 18352 11940 18358
rect 11888 18294 11940 18300
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11900 17882 11928 18294
rect 12256 18080 12308 18086
rect 12256 18022 12308 18028
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 12268 17678 12296 18022
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 10600 17604 10732 17610
rect 10652 17598 10732 17604
rect 10600 17546 10652 17552
rect 10704 17338 10732 17598
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10428 16182 10456 16730
rect 10876 16448 10928 16454
rect 10876 16390 10928 16396
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10048 16108 10100 16114
rect 10048 16050 10100 16056
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 10060 15570 10088 16050
rect 10048 15564 10100 15570
rect 10048 15506 10100 15512
rect 10060 15162 10088 15506
rect 10428 15434 10456 16118
rect 10888 16114 10916 16390
rect 10876 16108 10928 16114
rect 10876 16050 10928 16056
rect 11164 15978 11192 17546
rect 12912 17202 12940 18294
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12808 17128 12860 17134
rect 12808 17070 12860 17076
rect 12440 17060 12492 17066
rect 12440 17002 12492 17008
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11152 15972 11204 15978
rect 11152 15914 11204 15920
rect 10508 15904 10560 15910
rect 10508 15846 10560 15852
rect 10520 15570 10548 15846
rect 10508 15564 10560 15570
rect 10508 15506 10560 15512
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 11256 15162 11284 16050
rect 11532 15638 11560 16050
rect 11992 16046 12020 16526
rect 12452 16522 12480 17002
rect 12716 16992 12768 16998
rect 12716 16934 12768 16940
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11888 15972 11940 15978
rect 11888 15914 11940 15920
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11520 15632 11572 15638
rect 11520 15574 11572 15580
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9968 14618 9996 14826
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9324 12406 9444 12434
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8576 11280 8628 11286
rect 8576 11222 8628 11228
rect 7932 11144 7984 11150
rect 7932 11086 7984 11092
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 6644 10600 6696 10606
rect 6644 10542 6696 10548
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5632 9648 5684 9654
rect 5632 9590 5684 9596
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5460 8906 5488 9114
rect 5448 8900 5500 8906
rect 5448 8842 5500 8848
rect 5356 8832 5408 8838
rect 5540 8832 5592 8838
rect 5356 8774 5408 8780
rect 5460 8780 5540 8786
rect 5460 8774 5592 8780
rect 5264 8492 5316 8498
rect 5264 8434 5316 8440
rect 4908 7750 4936 7822
rect 5184 7806 5304 7834
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4540 6956 4660 6984
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4448 6322 4476 6802
rect 4540 6730 4568 6956
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4540 6458 4568 6666
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4632 6338 4660 6598
rect 4724 6440 4752 7142
rect 4816 6730 4844 7346
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4724 6412 4936 6440
rect 4436 6316 4488 6322
rect 4632 6310 4752 6338
rect 4436 6258 4488 6264
rect 4448 6202 4476 6258
rect 4448 6174 4660 6202
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4706 4660 6174
rect 4724 5914 4752 6310
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4816 5846 4844 6190
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4908 5658 4936 6412
rect 5276 5914 5304 7806
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5368 5846 5396 8774
rect 5460 8758 5580 8774
rect 5460 8362 5488 8758
rect 5644 8514 5672 9590
rect 6012 9382 6040 9862
rect 6000 9376 6052 9382
rect 6000 9318 6052 9324
rect 5644 8486 5764 8514
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5644 7886 5672 8366
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5552 7478 5580 7822
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 7002 5488 7142
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5356 5840 5408 5846
rect 5356 5782 5408 5788
rect 4816 5642 4936 5658
rect 4816 5636 4948 5642
rect 4816 5630 4896 5636
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4540 4690 4660 4706
rect 4528 4684 4660 4690
rect 4580 4678 4660 4684
rect 4528 4626 4580 4632
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4448 4282 4476 4490
rect 4632 4282 4660 4678
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4724 4214 4752 4966
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4816 3942 4844 5630
rect 4896 5578 4948 5584
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5368 5234 5396 5782
rect 5552 5302 5580 7414
rect 5736 7274 5764 8486
rect 5908 8492 5960 8498
rect 6012 8480 6040 9318
rect 6104 8974 6132 9998
rect 6656 9722 6684 10542
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 7024 9654 7052 9862
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 6092 8968 6144 8974
rect 6092 8910 6144 8916
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6274 8936 6330 8945
rect 6092 8560 6144 8566
rect 6196 8537 6224 8910
rect 6274 8871 6276 8880
rect 6328 8871 6330 8880
rect 6276 8842 6328 8848
rect 6092 8502 6144 8508
rect 6182 8528 6238 8537
rect 5960 8452 6040 8480
rect 5908 8434 5960 8440
rect 5816 8288 5868 8294
rect 5816 8230 5868 8236
rect 5828 7546 5856 8230
rect 6104 7886 6132 8502
rect 6182 8463 6184 8472
rect 6236 8463 6238 8472
rect 6184 8434 6236 8440
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5724 7268 5776 7274
rect 5724 7210 5776 7216
rect 6196 7002 6224 8434
rect 6288 7886 6316 8842
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6472 8362 6500 8434
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6748 7546 6776 8434
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6840 7478 6868 7958
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6932 7410 6960 7754
rect 7116 7410 7144 10406
rect 7760 10266 7788 10610
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 7748 10260 7800 10266
rect 7748 10202 7800 10208
rect 8128 10062 8156 10406
rect 8680 10062 8708 11018
rect 8956 10674 8984 11494
rect 9140 11150 9168 11562
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9324 11218 9352 11494
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8668 10056 8720 10062
rect 8668 9998 8720 10004
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 8576 9988 8628 9994
rect 8576 9930 8628 9936
rect 7392 8974 7420 9930
rect 8024 9036 8076 9042
rect 8392 9036 8444 9042
rect 8076 8996 8156 9024
rect 8024 8978 8076 8984
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8900 7340 8906
rect 7288 8842 7340 8848
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 7208 8430 7236 8774
rect 7300 8498 7328 8842
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7208 7886 7236 8366
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7392 7818 7420 8910
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7852 7818 7880 8434
rect 7944 8090 7972 8434
rect 7932 8084 7984 8090
rect 7932 8026 7984 8032
rect 8036 7886 8064 8502
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8128 7868 8156 8996
rect 8392 8978 8444 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8312 8634 8340 8910
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8220 8022 8248 8366
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8404 7886 8432 8978
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8496 8090 8524 8434
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8208 7880 8260 7886
rect 8128 7840 8208 7868
rect 7380 7812 7432 7818
rect 7380 7754 7432 7760
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 7116 6866 7144 7346
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6932 6458 6960 6734
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5276 4146 5304 4966
rect 5264 4140 5316 4146
rect 5368 4128 5396 5170
rect 5552 4826 5580 5238
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5448 4140 5500 4146
rect 5368 4100 5448 4128
rect 5264 4082 5316 4088
rect 5448 4082 5500 4088
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4816 3670 4844 3878
rect 5552 3738 5580 4558
rect 5828 4214 5856 4558
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5920 3942 5948 4762
rect 6656 4554 6684 4762
rect 6840 4622 6868 6258
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 4804 3664 4856 3670
rect 4804 3606 4856 3612
rect 5736 3466 5764 3878
rect 6196 3670 6224 3878
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6380 3602 6408 4422
rect 6472 4146 6500 4422
rect 6460 4140 6512 4146
rect 6460 4082 6512 4088
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 6380 2582 6408 3538
rect 6564 3058 6592 4082
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6840 3738 6868 4014
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6932 3466 6960 6394
rect 7668 6322 7696 7278
rect 7852 7274 7880 7754
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 8128 6458 8156 7840
rect 8208 7822 8260 7828
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8588 6866 8616 9930
rect 8864 9178 8892 10474
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 9048 9042 9076 10610
rect 9140 9110 9168 11086
rect 9416 11082 9444 12406
rect 9600 11830 9628 14282
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9784 12986 9812 13194
rect 9876 13190 9904 14010
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9692 12306 9720 12922
rect 9876 12918 9904 13126
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9876 12238 9904 12854
rect 10152 12782 10180 13670
rect 10140 12776 10192 12782
rect 10140 12718 10192 12724
rect 10152 12238 10180 12718
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 10140 12232 10192 12238
rect 10140 12174 10192 12180
rect 9876 11880 9904 12174
rect 9876 11852 9996 11880
rect 9588 11824 9640 11830
rect 9588 11766 9640 11772
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9496 10464 9548 10470
rect 9496 10406 9548 10412
rect 9508 10266 9536 10406
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9232 8498 9260 8842
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 8944 8356 8996 8362
rect 8944 8298 8996 8304
rect 8956 7886 8984 8298
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 7886 9260 8230
rect 9324 8090 9352 8910
rect 9416 8634 9444 8910
rect 9508 8634 9536 8978
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9416 7886 9444 8434
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9036 7744 9088 7750
rect 9036 7686 9088 7692
rect 9048 7546 9076 7686
rect 9416 7546 9444 7822
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9600 7478 9628 11766
rect 9864 11756 9916 11762
rect 9864 11698 9916 11704
rect 9876 11150 9904 11698
rect 9968 11694 9996 11852
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 10810 10088 11086
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9692 9654 9720 10678
rect 10152 10606 10180 11698
rect 10244 11558 10272 14758
rect 10888 14482 10916 15098
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 10336 13734 10364 14282
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10428 14006 10456 14214
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10416 14000 10468 14006
rect 10416 13942 10468 13948
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10324 13728 10376 13734
rect 10324 13670 10376 13676
rect 10336 12850 10364 13670
rect 10324 12844 10376 12850
rect 10324 12786 10376 12792
rect 10520 12238 10548 13806
rect 10704 13802 10732 14010
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10704 13530 10732 13738
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10888 13394 10916 14418
rect 10980 13734 11008 15098
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10704 12442 10732 12854
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10888 11762 10916 13330
rect 11072 12782 11100 14894
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11164 12986 11192 13194
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11348 12238 11376 15030
rect 11532 14958 11560 15574
rect 11624 15502 11652 15846
rect 11900 15586 11928 15914
rect 11992 15706 12020 15982
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12728 15638 12756 16934
rect 12820 16658 12848 17070
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12912 16114 12940 17138
rect 13096 16998 13124 18362
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 12992 16448 13044 16454
rect 12992 16390 13044 16396
rect 13004 16250 13032 16390
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 13096 16114 13124 16934
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12440 15632 12492 15638
rect 11900 15558 12020 15586
rect 12440 15574 12492 15580
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 11992 15094 12020 15558
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11992 14958 12020 15030
rect 12452 14958 12480 15574
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11808 12986 11836 13194
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11992 12646 12020 14894
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12452 14618 12480 14758
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12544 14550 12572 14962
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 14006 12112 14214
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12084 13190 12112 13806
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12452 12986 12480 13806
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 11980 12640 12032 12646
rect 11980 12582 12032 12588
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10796 11354 10824 11630
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10690 10732 10950
rect 10876 10736 10928 10742
rect 10704 10684 10876 10690
rect 10704 10678 10928 10684
rect 10704 10674 10916 10678
rect 10692 10668 10916 10674
rect 10744 10662 10916 10668
rect 10692 10610 10744 10616
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10152 10266 10180 10542
rect 10140 10260 10192 10266
rect 10140 10202 10192 10208
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9784 9518 9812 10066
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9784 8566 9812 9454
rect 10152 9178 10180 9522
rect 10140 9172 10192 9178
rect 10140 9114 10192 9120
rect 10428 9024 10456 9590
rect 10704 9178 10732 10610
rect 10980 10470 11008 11086
rect 11244 11076 11296 11082
rect 11244 11018 11296 11024
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11164 10674 11192 10950
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 10968 10464 11020 10470
rect 10968 10406 11020 10412
rect 10980 9586 11008 10406
rect 11164 10266 11192 10610
rect 11152 10260 11204 10266
rect 11152 10202 11204 10208
rect 11256 10062 11284 11018
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 11164 9466 11192 9522
rect 10980 9438 11192 9466
rect 10980 9178 11008 9438
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10600 9036 10652 9042
rect 10428 8996 10600 9024
rect 10600 8978 10652 8984
rect 10140 8900 10192 8906
rect 10140 8842 10192 8848
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9692 7886 9720 8230
rect 9784 7954 9812 8502
rect 9876 8498 9904 8774
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9680 7880 9732 7886
rect 9732 7828 9812 7834
rect 9680 7822 9812 7828
rect 9692 7806 9812 7822
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7656 6316 7708 6322
rect 7708 6276 7788 6304
rect 7656 6258 7708 6264
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7300 5710 7328 6054
rect 7484 5846 7512 6054
rect 7760 5846 7788 6276
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7748 5840 7800 5846
rect 7748 5782 7800 5788
rect 7760 5710 7788 5782
rect 7288 5704 7340 5710
rect 7288 5646 7340 5652
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7944 5234 7972 6326
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 6089 8064 6122
rect 8022 6080 8078 6089
rect 8022 6015 8078 6024
rect 8220 5710 8248 6734
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 8482 6352 8538 6361
rect 8300 6316 8352 6322
rect 8352 6296 8482 6304
rect 8352 6287 8538 6296
rect 8352 6276 8524 6287
rect 8300 6258 8352 6264
rect 8208 5704 8260 5710
rect 8128 5664 8208 5692
rect 8128 5574 8156 5664
rect 8208 5646 8260 5652
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8392 5636 8444 5642
rect 8392 5578 8444 5584
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8312 5302 8340 5578
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 8404 5166 8432 5578
rect 8496 5574 8524 6276
rect 8772 6202 8800 6394
rect 8850 6352 8906 6361
rect 8850 6287 8852 6296
rect 8904 6287 8906 6296
rect 8944 6316 8996 6322
rect 8852 6258 8904 6264
rect 8944 6258 8996 6264
rect 8680 6174 8800 6202
rect 8852 6180 8904 6186
rect 8680 6118 8708 6174
rect 8852 6122 8904 6128
rect 8668 6112 8720 6118
rect 8760 6112 8812 6118
rect 8668 6054 8720 6060
rect 8758 6080 8760 6089
rect 8812 6080 8814 6089
rect 8758 6015 8814 6024
rect 8864 5778 8892 6122
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8220 3670 8248 4014
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 7024 2650 7052 3606
rect 8220 3466 8248 3606
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7116 2650 7144 2926
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 7208 2378 7236 3334
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 8036 2650 8064 3062
rect 8128 2854 8156 3402
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 8128 2446 8156 2790
rect 8496 2582 8524 5170
rect 8680 2650 8708 5510
rect 8772 5234 8800 5578
rect 8760 5228 8812 5234
rect 8760 5170 8812 5176
rect 8772 4622 8800 5170
rect 8760 4616 8812 4622
rect 8760 4558 8812 4564
rect 8772 4282 8800 4558
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8864 4162 8892 5714
rect 8956 5234 8984 6258
rect 9128 5908 9180 5914
rect 9128 5850 9180 5856
rect 9036 5840 9088 5846
rect 9036 5782 9088 5788
rect 9048 5234 9076 5782
rect 9140 5574 9168 5850
rect 9324 5710 9352 6394
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 9036 5228 9088 5234
rect 9088 5188 9168 5216
rect 9036 5170 9088 5176
rect 8772 4134 8892 4162
rect 8956 4604 8984 5170
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 9048 4826 9076 5034
rect 9036 4820 9088 4826
rect 9036 4762 9088 4768
rect 9140 4690 9168 5188
rect 9324 4826 9352 5646
rect 9416 5234 9444 7346
rect 9600 6730 9628 7414
rect 9588 6724 9640 6730
rect 9588 6666 9640 6672
rect 9784 6662 9812 7806
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9876 6798 9904 6870
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 6322 9812 6598
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5302 9536 5646
rect 9680 5636 9732 5642
rect 9680 5578 9732 5584
rect 9692 5522 9720 5578
rect 9600 5494 9720 5522
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9416 4758 9444 5170
rect 9600 5166 9628 5494
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9404 4752 9456 4758
rect 9404 4694 9456 4700
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9036 4616 9088 4622
rect 8956 4576 9036 4604
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8484 2576 8536 2582
rect 8484 2518 8536 2524
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 7760 800 7788 2314
rect 8404 800 8432 2382
rect 8772 2310 8800 4134
rect 8852 3528 8904 3534
rect 8956 3516 8984 4576
rect 9036 4558 9088 4564
rect 9416 4282 9444 4694
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 8904 3488 8984 3516
rect 8852 3470 8904 3476
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8864 3126 8892 3334
rect 8852 3120 8904 3126
rect 8852 3062 8904 3068
rect 8956 2990 8984 3488
rect 9232 2990 9260 4082
rect 9416 3670 9444 4218
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9404 3664 9456 3670
rect 9404 3606 9456 3612
rect 9416 3534 9444 3606
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9232 2854 9260 2926
rect 9416 2854 9444 3470
rect 9692 3466 9720 4082
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9784 2582 9812 6258
rect 9876 6186 9904 6734
rect 9968 6390 9996 8366
rect 10060 7886 10088 8366
rect 10152 8090 10180 8842
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10324 8424 10376 8430
rect 10324 8366 10376 8372
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 10060 6322 10088 6802
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 10048 6180 10100 6186
rect 10048 6122 10100 6128
rect 9876 5914 9904 6122
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9956 5704 10008 5710
rect 9956 5646 10008 5652
rect 9968 5302 9996 5646
rect 10060 5642 10088 6122
rect 10152 6118 10180 7822
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9968 4146 9996 5238
rect 10152 5234 10180 5782
rect 10244 5370 10272 6258
rect 10336 5710 10364 8366
rect 10520 7750 10548 8434
rect 10612 7750 10640 8978
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10508 7744 10560 7750
rect 10506 7712 10508 7721
rect 10600 7744 10652 7750
rect 10560 7712 10562 7721
rect 10600 7686 10652 7692
rect 10506 7647 10562 7656
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 6662 10456 6734
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10612 6186 10640 7686
rect 10796 6798 10824 8774
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10888 7546 10916 7890
rect 10980 7886 11008 9114
rect 11256 8974 11284 9998
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11348 8906 11376 12174
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 11830 11928 12038
rect 12544 11898 12572 13806
rect 12636 13326 12664 13942
rect 12728 13462 12756 15438
rect 13188 15434 13216 16390
rect 13280 16250 13308 19314
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13452 18420 13504 18426
rect 13452 18362 13504 18368
rect 13464 18290 13492 18362
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17202 13400 18022
rect 13360 17196 13412 17202
rect 13360 17138 13412 17144
rect 13372 16658 13400 17138
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13268 16244 13320 16250
rect 13320 16204 13400 16232
rect 13268 16186 13320 16192
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 12808 14816 12860 14822
rect 12808 14758 12860 14764
rect 12820 14346 12848 14758
rect 12808 14340 12860 14346
rect 12808 14282 12860 14288
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12820 13530 12848 13874
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11808 11354 11836 11766
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 12912 11286 12940 15302
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 13004 14006 13032 14214
rect 13188 14006 13216 15370
rect 13280 15162 13308 16050
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13280 14482 13308 15098
rect 13372 14600 13400 16204
rect 13464 16114 13492 18090
rect 13556 18086 13584 18566
rect 13740 18290 13768 18566
rect 13832 18290 13860 21406
rect 14186 21382 14242 22182
rect 14830 21382 14886 22182
rect 14200 19514 14228 21382
rect 14844 20738 14872 21382
rect 14832 20732 14884 20738
rect 14832 20674 14884 20680
rect 16856 20732 16908 20738
rect 16856 20674 16908 20680
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15948 19378 15976 19450
rect 16868 19378 16896 20674
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 15936 19372 15988 19378
rect 15936 19314 15988 19320
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 14200 18766 14228 19314
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14292 18766 14320 19178
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14832 19168 14884 19174
rect 14832 19110 14884 19116
rect 14188 18760 14240 18766
rect 14188 18702 14240 18708
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 14200 17678 14228 18702
rect 14292 18426 14320 18702
rect 14384 18426 14412 19110
rect 14844 18766 14872 19110
rect 15396 18970 15424 19246
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 14832 18760 14884 18766
rect 14832 18702 14884 18708
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 14372 18420 14424 18426
rect 14844 18408 14872 18702
rect 15292 18692 15344 18698
rect 15292 18634 15344 18640
rect 14372 18362 14424 18368
rect 14752 18380 14872 18408
rect 15016 18420 15068 18426
rect 14752 17762 14780 18380
rect 15016 18362 15068 18368
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14568 17734 14780 17762
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16794 13768 16934
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 14292 16590 14320 17478
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14384 16794 14412 17138
rect 14372 16788 14424 16794
rect 14372 16730 14424 16736
rect 14568 16658 14596 17734
rect 14844 17678 14872 18226
rect 14924 17808 14976 17814
rect 14924 17750 14976 17756
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14660 17292 14872 17320
rect 14660 17202 14688 17292
rect 14738 17232 14794 17241
rect 14648 17196 14700 17202
rect 14844 17202 14872 17292
rect 14738 17167 14740 17176
rect 14648 17138 14700 17144
rect 14792 17167 14794 17176
rect 14832 17196 14884 17202
rect 14740 17138 14792 17144
rect 14832 17138 14884 17144
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 14384 16182 14412 16390
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 13464 15502 13492 16050
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13452 15496 13504 15502
rect 13452 15438 13504 15444
rect 13556 15162 13584 15914
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13556 15026 13584 15098
rect 13544 15020 13596 15026
rect 13544 14962 13596 14968
rect 13452 14612 13504 14618
rect 13372 14572 13452 14600
rect 13452 14554 13504 14560
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 13372 13938 13400 14418
rect 13464 14414 13492 14554
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13452 13932 13504 13938
rect 13740 13920 13768 14282
rect 13504 13892 13768 13920
rect 13452 13874 13504 13880
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 12992 13728 13044 13734
rect 12992 13670 13044 13676
rect 13004 13326 13032 13670
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13096 13258 13124 13738
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13372 12850 13400 13874
rect 13820 13864 13872 13870
rect 13740 13812 13820 13818
rect 13740 13806 13872 13812
rect 13740 13790 13860 13806
rect 13740 13530 13768 13790
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13728 13524 13780 13530
rect 13728 13466 13780 13472
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13556 12986 13584 13262
rect 13740 13190 13768 13466
rect 13832 13326 13860 13670
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13832 12782 13860 13262
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 14016 11762 14044 12854
rect 14476 12442 14504 16050
rect 14568 15910 14596 16594
rect 14660 16232 14688 17138
rect 14936 16590 14964 17750
rect 15028 17610 15056 18362
rect 15304 18290 15332 18634
rect 15488 18358 15516 19246
rect 15948 18834 15976 19314
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16132 18902 16160 19178
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16120 18896 16172 18902
rect 16120 18838 16172 18844
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 16316 18766 16344 19110
rect 16500 18766 16528 19178
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15304 17542 15332 18226
rect 15488 17678 15516 18294
rect 15764 18290 15792 18566
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15568 18080 15620 18086
rect 15568 18022 15620 18028
rect 15580 17678 15608 18022
rect 15764 17746 15792 18226
rect 15936 18148 15988 18154
rect 15936 18090 15988 18096
rect 15844 17808 15896 17814
rect 15844 17750 15896 17756
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 15120 17218 15148 17274
rect 15028 17202 15148 17218
rect 15016 17196 15148 17202
rect 15068 17190 15148 17196
rect 15198 17232 15254 17241
rect 15198 17167 15254 17176
rect 15016 17138 15068 17144
rect 15028 16998 15056 17138
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14924 16584 14976 16590
rect 14976 16544 15056 16572
rect 14924 16526 14976 16532
rect 14740 16244 14792 16250
rect 14660 16204 14740 16232
rect 14740 16186 14792 16192
rect 14924 16108 14976 16114
rect 14924 16050 14976 16056
rect 14936 15910 14964 16050
rect 15028 16046 15056 16544
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 15212 15978 15240 17167
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15200 15972 15252 15978
rect 15200 15914 15252 15920
rect 14556 15904 14608 15910
rect 14556 15846 14608 15852
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14660 12306 14688 12650
rect 14740 12640 14792 12646
rect 14936 12628 14964 15846
rect 15304 15502 15332 16118
rect 15396 16114 15424 16934
rect 15488 16590 15516 17070
rect 15856 17066 15884 17750
rect 15948 17202 15976 18090
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15580 16590 15608 17002
rect 15856 16590 15884 17002
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15948 16182 15976 17138
rect 16212 16448 16264 16454
rect 16212 16390 16264 16396
rect 15936 16176 15988 16182
rect 15936 16118 15988 16124
rect 16224 16114 16252 16390
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 15384 16108 15436 16114
rect 15384 16050 15436 16056
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 15936 15904 15988 15910
rect 15936 15846 15988 15852
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15488 15094 15516 15506
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15120 13138 15148 13874
rect 15212 13258 15240 13874
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15120 13110 15240 13138
rect 15016 12912 15068 12918
rect 15212 12866 15240 13110
rect 15016 12854 15068 12860
rect 14792 12600 14964 12628
rect 14740 12582 14792 12588
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 15028 12238 15056 12854
rect 15120 12838 15240 12866
rect 15120 12374 15148 12838
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15212 12306 15240 12582
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 12900 11280 12952 11286
rect 12900 11222 12952 11228
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 11428 11076 11480 11082
rect 11428 11018 11480 11024
rect 11440 10810 11468 11018
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 12360 10674 12388 10950
rect 13188 10810 13216 11086
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13188 10674 13216 10746
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 13096 10198 13124 10406
rect 13084 10192 13136 10198
rect 13084 10134 13136 10140
rect 13280 10062 13308 11630
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13820 11552 13872 11558
rect 13820 11494 13872 11500
rect 13912 11552 13964 11558
rect 13912 11494 13964 11500
rect 13556 11150 13584 11494
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13372 10470 13400 11086
rect 13464 10810 13492 11086
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13832 10606 13860 11494
rect 13924 11218 13952 11494
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 14016 11150 14044 11698
rect 14108 11354 14136 11698
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 15304 11150 15332 14758
rect 15396 12434 15424 14962
rect 15488 14890 15516 15030
rect 15476 14884 15528 14890
rect 15476 14826 15528 14832
rect 15764 14618 15792 15438
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15488 12850 15516 14554
rect 15856 14414 15884 14758
rect 15948 14482 15976 15846
rect 16224 15638 16252 16050
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14482 16436 14758
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16132 12986 16160 13874
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15672 12646 15700 12922
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15936 12436 15988 12442
rect 15396 12406 15516 12434
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 14004 11144 14056 11150
rect 14004 11086 14056 11092
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14660 10674 14688 10746
rect 15016 10736 15068 10742
rect 15014 10704 15016 10713
rect 15200 10736 15252 10742
rect 15068 10704 15070 10713
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14648 10668 14700 10674
rect 15200 10678 15252 10684
rect 15014 10639 15070 10648
rect 14648 10610 14700 10616
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13372 10266 13400 10406
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 12992 10056 13044 10062
rect 12992 9998 13044 10004
rect 13268 10056 13320 10062
rect 13268 9998 13320 10004
rect 12256 9648 12308 9654
rect 12256 9590 12308 9596
rect 12268 9178 12296 9590
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 10968 7880 11020 7886
rect 10968 7822 11020 7828
rect 10980 7546 11008 7822
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6458 10824 6734
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5710 10548 6054
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10232 5364 10284 5370
rect 10232 5306 10284 5312
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10140 4004 10192 4010
rect 10140 3946 10192 3952
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10152 3738 10180 3946
rect 10140 3732 10192 3738
rect 10140 3674 10192 3680
rect 10428 3602 10456 3946
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10152 3194 10180 3470
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10520 3126 10548 4150
rect 10612 3942 10640 6122
rect 10704 5234 10732 6258
rect 10796 6254 10824 6394
rect 10888 6254 10916 7482
rect 11532 6984 11560 8502
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11624 8090 11652 8230
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 12072 7948 12124 7954
rect 12072 7890 12124 7896
rect 12084 7478 12112 7890
rect 12176 7478 12204 8910
rect 13004 8634 13032 9998
rect 13648 9722 13676 10406
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13912 9716 13964 9722
rect 13912 9658 13964 9664
rect 13924 9586 13952 9658
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 13820 9444 13872 9450
rect 13820 9386 13872 9392
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12256 7812 12308 7818
rect 12256 7754 12308 7760
rect 12268 7546 12296 7754
rect 12360 7750 12388 8298
rect 13280 7750 13308 8366
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11612 6996 11664 7002
rect 11532 6956 11612 6984
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 6361 11192 6598
rect 11150 6352 11206 6361
rect 11532 6322 11560 6956
rect 11612 6938 11664 6944
rect 11612 6860 11664 6866
rect 11612 6802 11664 6808
rect 11624 6458 11652 6802
rect 11808 6662 11836 7346
rect 11992 7274 12020 7346
rect 11980 7268 12032 7274
rect 11980 7210 12032 7216
rect 11992 6712 12020 7210
rect 12084 6984 12112 7414
rect 12176 7206 12204 7414
rect 12360 7342 12388 7686
rect 13280 7478 13308 7686
rect 13464 7546 13492 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13268 7472 13320 7478
rect 13268 7414 13320 7420
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12164 6996 12216 7002
rect 12084 6956 12164 6984
rect 12164 6938 12216 6944
rect 12072 6724 12124 6730
rect 11992 6684 12072 6712
rect 12072 6666 12124 6672
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11150 6287 11152 6296
rect 11204 6287 11206 6296
rect 11520 6316 11572 6322
rect 11152 6258 11204 6264
rect 11520 6258 11572 6264
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5914 11008 6054
rect 11992 5914 12020 6326
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 10876 5772 10928 5778
rect 10796 5732 10876 5760
rect 10796 5574 10824 5732
rect 10876 5714 10928 5720
rect 12084 5710 12112 6666
rect 12636 6662 12664 7142
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12360 5778 12388 6598
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10876 5568 10928 5574
rect 10876 5510 10928 5516
rect 12164 5568 12216 5574
rect 12164 5510 12216 5516
rect 10888 5370 10916 5510
rect 10876 5364 10928 5370
rect 10876 5306 10928 5312
rect 12176 5302 12204 5510
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10416 3120 10468 3126
rect 10414 3088 10416 3097
rect 10508 3120 10560 3126
rect 10468 3088 10470 3097
rect 10508 3062 10560 3068
rect 10414 3023 10470 3032
rect 10612 2854 10640 3878
rect 10704 3058 10732 4082
rect 11072 3398 11100 4150
rect 12176 4146 12204 5238
rect 12268 5234 12296 5578
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12360 4622 12388 5714
rect 12544 5234 12572 6190
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12348 4616 12400 4622
rect 12268 4576 12348 4604
rect 12268 4282 12296 4576
rect 12348 4558 12400 4564
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 12360 4146 12388 4422
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12544 4128 12572 5170
rect 12636 4622 12664 6598
rect 12728 5710 12756 6938
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 6390 13492 6598
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13556 5710 13584 8842
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 7750 13768 8434
rect 13832 8362 13860 9386
rect 14016 8634 14044 10610
rect 14660 10062 14688 10610
rect 15212 10554 15240 10678
rect 15396 10674 15424 11494
rect 15384 10668 15436 10674
rect 15384 10610 15436 10616
rect 15120 10526 15240 10554
rect 15384 10532 15436 10538
rect 15120 10130 15148 10526
rect 15384 10474 15436 10480
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15212 10062 15240 10406
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14648 10056 14700 10062
rect 15200 10056 15252 10062
rect 14648 9998 14700 10004
rect 15106 10024 15162 10033
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 13912 8492 13964 8498
rect 13912 8434 13964 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13924 8022 13952 8434
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 13912 8016 13964 8022
rect 13912 7958 13964 7964
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 14016 7546 14044 8366
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13832 7274 13860 7346
rect 14108 7274 14136 8502
rect 14200 8090 14228 9998
rect 14292 9518 14320 9998
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 14384 9586 14412 9862
rect 14660 9722 14688 9998
rect 15200 9998 15252 10004
rect 15106 9959 15162 9968
rect 15120 9926 15148 9959
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15200 9920 15252 9926
rect 15200 9862 15252 9868
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 14384 8498 14412 9522
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 15108 8016 15160 8022
rect 15028 7976 15108 8004
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14384 7410 14412 7890
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14832 7880 14884 7886
rect 14832 7822 14884 7828
rect 14476 7478 14504 7822
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14568 7410 14596 7754
rect 14844 7410 14872 7822
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14936 7410 14964 7686
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 13832 6458 13860 7210
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 14844 6322 14872 7346
rect 15028 7206 15056 7976
rect 15108 7958 15160 7964
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15120 7206 15148 7482
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15028 6662 15056 7142
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 14832 6316 14884 6322
rect 14832 6258 14884 6264
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14568 5710 14596 6190
rect 12716 5704 12768 5710
rect 12716 5646 12768 5652
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13648 4826 13676 5238
rect 14476 5030 14504 5510
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 13820 4208 13872 4214
rect 13820 4150 13872 4156
rect 12624 4140 12676 4146
rect 12544 4100 12624 4128
rect 11716 3602 11744 4082
rect 11900 3738 11928 4082
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 11072 3058 11100 3334
rect 11532 3126 11560 3470
rect 12084 3398 12112 4014
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 11520 3120 11572 3126
rect 11150 3088 11206 3097
rect 10692 3052 10744 3058
rect 10692 2994 10744 3000
rect 11060 3052 11112 3058
rect 11520 3062 11572 3068
rect 12084 3058 12112 3334
rect 12360 3126 12388 3674
rect 12544 3194 12572 4100
rect 12624 4082 12676 4088
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12636 3534 12664 3946
rect 13832 3738 13860 4150
rect 14568 3942 14596 5646
rect 14648 5636 14700 5642
rect 14648 5578 14700 5584
rect 14660 5302 14688 5578
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14844 5234 14872 6258
rect 15120 6254 15148 7142
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15212 5914 15240 9862
rect 15304 9722 15332 10066
rect 15396 10010 15424 10474
rect 15488 10266 15516 12406
rect 15936 12378 15988 12384
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15672 12186 15700 12242
rect 15948 12238 15976 12378
rect 16040 12238 16068 12650
rect 16132 12442 16160 12718
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 15936 12232 15988 12238
rect 15672 12158 15792 12186
rect 15936 12174 15988 12180
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15764 12102 15792 12158
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15764 11762 15792 12038
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15764 11354 15792 11698
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 15660 10668 15712 10674
rect 15580 10628 15660 10656
rect 15476 10260 15528 10266
rect 15476 10202 15528 10208
rect 15580 10010 15608 10628
rect 15660 10610 15712 10616
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15396 9994 15608 10010
rect 15384 9988 15608 9994
rect 15436 9982 15608 9988
rect 15384 9930 15436 9936
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15580 9654 15608 9982
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15672 9586 15700 10474
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9722 15792 9998
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15488 9450 15516 9522
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15488 9178 15516 9386
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15488 7818 15516 8434
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15476 7812 15528 7818
rect 15476 7754 15528 7760
rect 15488 7274 15516 7754
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 15384 7200 15436 7206
rect 15384 7142 15436 7148
rect 15396 6322 15424 7142
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15212 5234 15240 5714
rect 15396 5710 15424 6258
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15488 5302 15516 6326
rect 15580 6254 15608 7822
rect 15856 6610 15884 11086
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10742 15976 10950
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15948 10146 15976 10678
rect 16040 10554 16068 11494
rect 16120 11008 16172 11014
rect 16120 10950 16172 10956
rect 16132 10674 16160 10950
rect 16120 10668 16172 10674
rect 16120 10610 16172 10616
rect 16040 10526 16160 10554
rect 15948 10118 16068 10146
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15672 6582 15884 6610
rect 15568 6248 15620 6254
rect 15568 6190 15620 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5914 15608 6054
rect 15568 5908 15620 5914
rect 15568 5850 15620 5856
rect 15476 5296 15528 5302
rect 15476 5238 15528 5244
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 11150 3023 11152 3032
rect 11060 2994 11112 3000
rect 11204 3023 11206 3032
rect 12072 3052 12124 3058
rect 11152 2994 11204 3000
rect 12072 2994 12124 3000
rect 13556 2854 13584 3334
rect 10600 2848 10652 2854
rect 10600 2790 10652 2796
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 13648 2446 13676 3470
rect 14844 3466 14872 5170
rect 15580 5030 15608 5850
rect 15672 5778 15700 6582
rect 15948 6458 15976 9998
rect 16040 9926 16068 10118
rect 16028 9920 16080 9926
rect 16028 9862 16080 9868
rect 16040 9518 16068 9862
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16132 7886 16160 10526
rect 16224 10266 16252 14350
rect 16592 14346 16620 15370
rect 16684 15026 16712 16186
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17316 15496 17368 15502
rect 17316 15438 17368 15444
rect 16672 15020 16724 15026
rect 16672 14962 16724 14968
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 16672 14884 16724 14890
rect 16672 14826 16724 14832
rect 16684 14618 16712 14826
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16684 14362 16712 14554
rect 17052 14414 17080 14962
rect 17236 14618 17264 14962
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17040 14408 17092 14414
rect 16580 14340 16632 14346
rect 16684 14334 16804 14362
rect 17040 14350 17092 14356
rect 16580 14282 16632 14288
rect 16672 14272 16724 14278
rect 16672 14214 16724 14220
rect 16684 14074 16712 14214
rect 16776 14074 16804 14334
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 17052 13870 17080 14350
rect 17328 14346 17356 15438
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17604 15162 17632 15302
rect 17788 15162 17816 15642
rect 17960 15428 18012 15434
rect 17960 15370 18012 15376
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17776 15156 17828 15162
rect 17776 15098 17828 15104
rect 17408 15088 17460 15094
rect 17408 15030 17460 15036
rect 17420 14618 17448 15030
rect 17972 14890 18000 15370
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18328 15020 18380 15026
rect 18328 14962 18380 14968
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 17960 14884 18012 14890
rect 17960 14826 18012 14832
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17972 14550 18000 14826
rect 17960 14544 18012 14550
rect 17960 14486 18012 14492
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17328 13530 17356 14282
rect 17788 13870 17816 14418
rect 18064 14362 18092 14962
rect 18340 14618 18368 14962
rect 18328 14612 18380 14618
rect 18328 14554 18380 14560
rect 18236 14408 18288 14414
rect 17972 14346 18092 14362
rect 17960 14340 18092 14346
rect 18012 14334 18092 14340
rect 18234 14376 18236 14385
rect 18288 14376 18290 14385
rect 18234 14311 18290 14320
rect 17960 14282 18012 14288
rect 17868 14272 17920 14278
rect 17868 14214 17920 14220
rect 17880 13938 17908 14214
rect 18340 14074 18368 14554
rect 18432 14482 18460 14962
rect 18420 14476 18472 14482
rect 18420 14418 18472 14424
rect 18432 14074 18460 14418
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17776 13864 17828 13870
rect 17776 13806 17828 13812
rect 17684 13796 17736 13802
rect 17684 13738 17736 13744
rect 17500 13728 17552 13734
rect 17500 13670 17552 13676
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 16580 13388 16632 13394
rect 16580 13330 16632 13336
rect 16592 12986 16620 13330
rect 17512 13326 17540 13670
rect 17696 13394 17724 13738
rect 17880 13734 17908 13874
rect 17868 13728 17920 13734
rect 18524 13705 18552 14350
rect 17868 13670 17920 13676
rect 18510 13696 18566 13705
rect 18510 13631 18566 13640
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16592 12782 16620 12922
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 17408 12844 17460 12850
rect 17408 12786 17460 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16776 12170 16804 12786
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 17052 12442 17080 12718
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17420 12238 17448 12786
rect 17512 12628 17540 12854
rect 18432 12850 18460 13126
rect 18524 13025 18552 13262
rect 18510 13016 18566 13025
rect 18510 12951 18566 12960
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 17592 12640 17644 12646
rect 17512 12600 17592 12628
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16776 11558 16804 12106
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16316 10742 16344 11222
rect 16868 11082 16896 11698
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16960 11082 16988 11630
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16408 10674 16436 11018
rect 16868 10810 16896 11018
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 17236 10742 17264 10950
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 17224 10736 17276 10742
rect 17224 10678 17276 10684
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 10266 16344 10406
rect 16408 10266 16436 10610
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 16396 10260 16448 10266
rect 16396 10202 16448 10208
rect 16316 9382 16344 10202
rect 16500 10198 16528 10678
rect 17236 10606 17264 10678
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17144 10470 17172 10542
rect 17132 10464 17184 10470
rect 17132 10406 17184 10412
rect 16488 10192 16540 10198
rect 16488 10134 16540 10140
rect 16396 10056 16448 10062
rect 17144 10033 17172 10406
rect 17236 10062 17264 10542
rect 17328 10062 17356 10678
rect 17224 10056 17276 10062
rect 16396 9998 16448 10004
rect 17130 10024 17186 10033
rect 16408 9926 16436 9998
rect 17224 9998 17276 10004
rect 17316 10056 17368 10062
rect 17316 9998 17368 10004
rect 17130 9959 17186 9968
rect 17144 9926 17172 9959
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17224 9648 17276 9654
rect 17224 9590 17276 9596
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 17236 9042 17264 9590
rect 17328 9178 17356 9998
rect 17420 9450 17448 12174
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17224 9036 17276 9042
rect 17276 8996 17356 9024
rect 17224 8978 17276 8984
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16028 7880 16080 7886
rect 16028 7822 16080 7828
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16040 7732 16068 7822
rect 16224 7750 16252 8774
rect 16868 8634 16896 8910
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16580 8016 16632 8022
rect 16632 7964 16712 7970
rect 16580 7958 16712 7964
rect 16592 7942 16712 7958
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16580 7880 16632 7886
rect 16580 7822 16632 7828
rect 16316 7750 16344 7822
rect 16212 7744 16264 7750
rect 16040 7704 16160 7732
rect 16132 7274 16160 7704
rect 16210 7712 16212 7721
rect 16304 7744 16356 7750
rect 16264 7712 16266 7721
rect 16304 7686 16356 7692
rect 16210 7647 16266 7656
rect 16120 7268 16172 7274
rect 16120 7210 16172 7216
rect 16592 6866 16620 7822
rect 16684 7410 16712 7942
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16776 7410 16804 7686
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16764 7404 16816 7410
rect 16764 7346 16816 7352
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16684 6798 16712 7346
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 16224 6322 16252 6598
rect 15844 6316 15896 6322
rect 16212 6316 16264 6322
rect 15844 6258 15896 6264
rect 16132 6276 16212 6304
rect 15856 6118 15884 6258
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15844 6112 15896 6118
rect 15844 6054 15896 6060
rect 15764 5778 15792 6054
rect 15660 5772 15712 5778
rect 15660 5714 15712 5720
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5370 15792 5714
rect 15936 5704 15988 5710
rect 16040 5692 16068 6122
rect 16132 5710 16160 6276
rect 16212 6258 16264 6264
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 15988 5664 16068 5692
rect 15936 5646 15988 5652
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 16040 5234 16068 5664
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16132 5370 16160 5646
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16028 5228 16080 5234
rect 16028 5170 16080 5176
rect 16224 5166 16252 5850
rect 16212 5160 16264 5166
rect 16212 5102 16264 5108
rect 16316 5098 16344 6258
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16408 5846 16436 6190
rect 16396 5840 16448 5846
rect 16396 5782 16448 5788
rect 16500 5370 16528 6258
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16592 5710 16620 6190
rect 16776 6118 16804 6870
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 16776 5710 16804 6054
rect 17052 5914 17080 8434
rect 17236 7954 17264 8774
rect 17328 8362 17356 8996
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17316 8356 17368 8362
rect 17316 8298 17368 8304
rect 17420 8294 17448 8910
rect 17512 8498 17540 12600
rect 17592 12582 17644 12588
rect 17684 12640 17736 12646
rect 17684 12582 17736 12588
rect 17696 12238 17724 12582
rect 18510 12336 18566 12345
rect 18510 12271 18566 12280
rect 18524 12238 18552 12271
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17590 10704 17646 10713
rect 17590 10639 17646 10648
rect 17604 10606 17632 10639
rect 17592 10600 17644 10606
rect 17592 10542 17644 10548
rect 17604 10198 17632 10542
rect 17592 10192 17644 10198
rect 17592 10134 17644 10140
rect 17972 10130 18000 10950
rect 18248 10305 18276 11086
rect 18328 11008 18380 11014
rect 18524 10985 18552 11086
rect 18328 10950 18380 10956
rect 18510 10976 18566 10985
rect 18340 10674 18368 10950
rect 18510 10911 18566 10920
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18234 10296 18290 10305
rect 18340 10266 18368 10610
rect 18234 10231 18290 10240
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 18340 10146 18368 10202
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 18248 10118 18368 10146
rect 17972 9586 18000 10066
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 18064 9178 18092 9454
rect 18248 9382 18276 10118
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18340 9722 18368 9998
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18340 9042 18368 9658
rect 18510 9616 18566 9625
rect 18510 9551 18512 9560
rect 18564 9551 18566 9560
rect 18512 9522 18564 9528
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 18236 8968 18288 8974
rect 18236 8910 18288 8916
rect 18418 8936 18474 8945
rect 17684 8900 17736 8906
rect 17684 8842 17736 8848
rect 18052 8900 18104 8906
rect 18052 8842 18104 8848
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 8022 17448 8230
rect 17512 8022 17540 8434
rect 17408 8016 17460 8022
rect 17408 7958 17460 7964
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7410 17172 7822
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17144 7274 17172 7346
rect 17236 7274 17264 7890
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 17224 7268 17276 7274
rect 17224 7210 17276 7216
rect 17316 7200 17368 7206
rect 17316 7142 17368 7148
rect 17222 6896 17278 6905
rect 17222 6831 17278 6840
rect 17236 6798 17264 6831
rect 17328 6798 17356 7142
rect 17224 6792 17276 6798
rect 17224 6734 17276 6740
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17316 6656 17368 6662
rect 17316 6598 17368 6604
rect 17222 6352 17278 6361
rect 17222 6287 17278 6296
rect 17236 6254 17264 6287
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17328 6118 17356 6598
rect 17420 6322 17448 7958
rect 17500 7880 17552 7886
rect 17604 7868 17632 8774
rect 17696 8634 17724 8842
rect 17684 8628 17736 8634
rect 17684 8570 17736 8576
rect 18064 8498 18092 8842
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18248 8430 18276 8910
rect 18418 8871 18474 8880
rect 18432 8566 18460 8871
rect 18524 8634 18552 9114
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18420 8560 18472 8566
rect 18420 8502 18472 8508
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17880 7954 17908 8230
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17552 7840 17632 7868
rect 17500 7822 17552 7828
rect 17512 7478 17540 7822
rect 17972 7546 18000 8298
rect 18248 8294 18276 8366
rect 18236 8288 18288 8294
rect 18236 8230 18288 8236
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18602 8256 18658 8265
rect 18432 7886 18460 8230
rect 18602 8191 18658 8200
rect 18420 7880 18472 7886
rect 18420 7822 18472 7828
rect 18050 7576 18106 7585
rect 17960 7540 18012 7546
rect 18050 7511 18106 7520
rect 17960 7482 18012 7488
rect 17500 7472 17552 7478
rect 17500 7414 17552 7420
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17408 6316 17460 6322
rect 17408 6258 17460 6264
rect 17512 6254 17540 7414
rect 17604 7002 17632 7414
rect 17972 7274 18000 7482
rect 18064 7342 18092 7511
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17960 7268 18012 7274
rect 17960 7210 18012 7216
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 18432 6798 18460 7822
rect 18420 6792 18472 6798
rect 18420 6734 18472 6740
rect 17500 6248 17552 6254
rect 18512 6248 18564 6254
rect 17500 6190 17552 6196
rect 18510 6216 18512 6225
rect 18564 6216 18566 6225
rect 18510 6151 18566 6160
rect 17316 6112 17368 6118
rect 17316 6054 17368 6060
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17328 5710 17356 6054
rect 18616 5710 18644 8191
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 16764 5704 16816 5710
rect 16764 5646 16816 5652
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 18604 5704 18656 5710
rect 18604 5646 18656 5652
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16868 5302 16896 5578
rect 17132 5568 17184 5574
rect 17132 5510 17184 5516
rect 16856 5296 16908 5302
rect 16856 5238 16908 5244
rect 17144 5234 17172 5510
rect 17132 5228 17184 5234
rect 17132 5170 17184 5176
rect 16304 5092 16356 5098
rect 16304 5034 16356 5040
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 3194 14872 3402
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 14016 2650 14044 3062
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 9048 800 9076 2314
rect 9692 800 9720 2382
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
<< via2 >>
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 1398 17720 1454 17776
rect 846 15816 902 15872
rect 846 14864 902 14920
rect 846 14456 902 14512
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 846 13132 848 13152
rect 848 13132 900 13152
rect 900 13132 902 13152
rect 846 13096 902 13132
rect 846 12180 848 12200
rect 848 12180 900 12200
rect 900 12180 902 12200
rect 846 12144 902 12180
rect 846 11756 902 11792
rect 846 11736 848 11756
rect 848 11736 900 11756
rect 900 11736 902 11756
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 846 10376 902 10432
rect 1398 9560 1454 9616
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 8022 18264 8078 18320
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 846 9016 902 9072
rect 2134 8916 2136 8936
rect 2136 8916 2188 8936
rect 2188 8916 2190 8936
rect 2134 8880 2190 8916
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1398 8200 1454 8256
rect 846 7656 902 7712
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3790 8492 3846 8528
rect 3790 8472 3792 8492
rect 3792 8472 3844 8492
rect 3844 8472 3846 8492
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 6274 8900 6330 8936
rect 6274 8880 6276 8900
rect 6276 8880 6328 8900
rect 6328 8880 6330 8900
rect 6182 8492 6238 8528
rect 6182 8472 6184 8492
rect 6184 8472 6236 8492
rect 6236 8472 6238 8492
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8022 6024 8078 6080
rect 8482 6296 8538 6352
rect 8850 6316 8906 6352
rect 8850 6296 8852 6316
rect 8852 6296 8904 6316
rect 8904 6296 8906 6316
rect 8758 6060 8760 6080
rect 8760 6060 8812 6080
rect 8812 6060 8814 6080
rect 8758 6024 8814 6060
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 10506 7692 10508 7712
rect 10508 7692 10560 7712
rect 10560 7692 10562 7712
rect 10506 7656 10562 7692
rect 14738 17196 14794 17232
rect 14738 17176 14740 17196
rect 14740 17176 14792 17196
rect 14792 17176 14794 17196
rect 15198 17176 15254 17232
rect 15014 10684 15016 10704
rect 15016 10684 15068 10704
rect 15068 10684 15070 10704
rect 15014 10648 15070 10684
rect 11150 6316 11206 6352
rect 11150 6296 11152 6316
rect 11152 6296 11204 6316
rect 11204 6296 11206 6316
rect 10414 3068 10416 3088
rect 10416 3068 10468 3088
rect 10468 3068 10470 3088
rect 10414 3032 10470 3068
rect 15106 9968 15162 10024
rect 11150 3052 11206 3088
rect 11150 3032 11152 3052
rect 11152 3032 11204 3052
rect 11204 3032 11206 3052
rect 18234 14356 18236 14376
rect 18236 14356 18288 14376
rect 18288 14356 18290 14376
rect 18234 14320 18290 14356
rect 18510 13640 18566 13696
rect 18510 12960 18566 13016
rect 17130 9968 17186 10024
rect 16210 7692 16212 7712
rect 16212 7692 16264 7712
rect 16264 7692 16266 7712
rect 16210 7656 16266 7692
rect 18510 12280 18566 12336
rect 17590 10648 17646 10704
rect 18510 10920 18566 10976
rect 18234 10240 18290 10296
rect 18510 9580 18566 9616
rect 18510 9560 18512 9580
rect 18512 9560 18564 9580
rect 18564 9560 18566 9580
rect 17222 6840 17278 6896
rect 17222 6296 17278 6352
rect 18418 8880 18474 8936
rect 18602 8200 18658 8256
rect 18050 7520 18106 7576
rect 18510 6196 18512 6216
rect 18512 6196 18564 6216
rect 18564 6196 18566 6216
rect 18510 6160 18566 6196
<< metal3 >>
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 0 18458 800 18488
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 0 18398 2790 18458
rect 0 18368 800 18398
rect 2730 18322 2790 18398
rect 8017 18322 8083 18325
rect 2730 18320 8083 18322
rect 2730 18264 8022 18320
rect 8078 18264 8083 18320
rect 2730 18262 8083 18264
rect 8017 18259 8083 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 14733 17234 14799 17237
rect 15193 17234 15259 17237
rect 14733 17232 15259 17234
rect 14733 17176 14738 17232
rect 14794 17176 15198 17232
rect 15254 17176 15259 17232
rect 14733 17174 15259 17176
rect 14733 17171 14799 17174
rect 15193 17171 15259 17174
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 841 15874 907 15877
rect 798 15872 907 15874
rect 798 15816 846 15872
rect 902 15816 907 15872
rect 798 15811 907 15816
rect 798 15768 858 15811
rect 0 15678 858 15768
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 0 15648 800 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 0 15058 800 15088
rect 0 14968 858 15058
rect 798 14925 858 14968
rect 798 14920 907 14925
rect 798 14864 846 14920
rect 902 14864 907 14920
rect 798 14862 907 14864
rect 841 14859 907 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 18229 14378 18295 14381
rect 19238 14378 20038 14408
rect 18229 14376 20038 14378
rect 18229 14320 18234 14376
rect 18290 14320 20038 14376
rect 18229 14318 20038 14320
rect 0 14288 800 14318
rect 18229 14315 18295 14318
rect 19238 14288 20038 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 18505 13698 18571 13701
rect 19238 13698 20038 13728
rect 18505 13696 20038 13698
rect 18505 13640 18510 13696
rect 18566 13640 20038 13696
rect 18505 13638 20038 13640
rect 18505 13635 18571 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 19238 13608 20038 13638
rect 4210 13567 4526 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 18505 13018 18571 13021
rect 19238 13018 20038 13048
rect 18505 13016 20038 13018
rect 18505 12960 18510 13016
rect 18566 12960 20038 13016
rect 18505 12958 20038 12960
rect 0 12928 800 12958
rect 18505 12955 18571 12958
rect 19238 12928 20038 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 0 12338 800 12368
rect 18505 12338 18571 12341
rect 19238 12338 20038 12368
rect 0 12248 858 12338
rect 18505 12336 20038 12338
rect 18505 12280 18510 12336
rect 18566 12280 20038 12336
rect 18505 12278 20038 12280
rect 18505 12275 18571 12278
rect 19238 12248 20038 12278
rect 798 12205 858 12248
rect 798 12200 907 12205
rect 798 12144 846 12200
rect 902 12144 907 12200
rect 798 12142 907 12144
rect 841 12139 907 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 0 11568 800 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 18505 10978 18571 10981
rect 19238 10978 20038 11008
rect 18505 10976 20038 10978
rect 18505 10920 18510 10976
rect 18566 10920 20038 10976
rect 18505 10918 20038 10920
rect 18505 10915 18571 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 19238 10888 20038 10918
rect 4870 10847 5186 10848
rect 15009 10706 15075 10709
rect 17585 10706 17651 10709
rect 15009 10704 17651 10706
rect 15009 10648 15014 10704
rect 15070 10648 17590 10704
rect 17646 10648 17651 10704
rect 15009 10646 17651 10648
rect 15009 10643 15075 10646
rect 17585 10643 17651 10646
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 18229 10298 18295 10301
rect 19238 10298 20038 10328
rect 18229 10296 20038 10298
rect 18229 10240 18234 10296
rect 18290 10240 20038 10296
rect 18229 10238 20038 10240
rect 0 10208 800 10238
rect 18229 10235 18295 10238
rect 19238 10208 20038 10238
rect 15101 10026 15167 10029
rect 17125 10026 17191 10029
rect 15101 10024 17191 10026
rect 15101 9968 15106 10024
rect 15162 9968 17130 10024
rect 17186 9968 17191 10024
rect 15101 9966 17191 9968
rect 15101 9963 15167 9966
rect 17125 9963 17191 9966
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 18505 9618 18571 9621
rect 19238 9618 20038 9648
rect 18505 9616 20038 9618
rect 18505 9560 18510 9616
rect 18566 9560 20038 9616
rect 18505 9558 20038 9560
rect 18505 9555 18571 9558
rect 19238 9528 20038 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 2129 8938 2195 8941
rect 6269 8938 6335 8941
rect 2129 8936 6335 8938
rect 2129 8880 2134 8936
rect 2190 8880 6274 8936
rect 6330 8880 6335 8936
rect 2129 8878 6335 8880
rect 0 8848 800 8878
rect 2129 8875 2195 8878
rect 6269 8875 6335 8878
rect 18413 8938 18479 8941
rect 19238 8938 20038 8968
rect 18413 8936 20038 8938
rect 18413 8880 18418 8936
rect 18474 8880 20038 8936
rect 18413 8878 20038 8880
rect 18413 8875 18479 8878
rect 19238 8848 20038 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 3785 8530 3851 8533
rect 6177 8530 6243 8533
rect 3785 8528 6243 8530
rect 3785 8472 3790 8528
rect 3846 8472 6182 8528
rect 6238 8472 6243 8528
rect 3785 8470 6243 8472
rect 3785 8467 3851 8470
rect 6177 8467 6243 8470
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 18597 8258 18663 8261
rect 19238 8258 20038 8288
rect 18597 8256 20038 8258
rect 18597 8200 18602 8256
rect 18658 8200 20038 8256
rect 18597 8198 20038 8200
rect 18597 8195 18663 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 19238 8168 20038 8198
rect 4210 8127 4526 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 10501 7714 10567 7717
rect 16205 7714 16271 7717
rect 10501 7712 16271 7714
rect 10501 7656 10506 7712
rect 10562 7656 16210 7712
rect 16266 7656 16271 7712
rect 10501 7654 16271 7656
rect 10501 7651 10567 7654
rect 16205 7651 16271 7654
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 18045 7578 18111 7581
rect 19238 7578 20038 7608
rect 18045 7576 20038 7578
rect 18045 7520 18050 7576
rect 18106 7520 20038 7576
rect 18045 7518 20038 7520
rect 0 7488 800 7518
rect 18045 7515 18111 7518
rect 19238 7488 20038 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 17217 6898 17283 6901
rect 19238 6898 20038 6928
rect 17217 6896 20038 6898
rect 17217 6840 17222 6896
rect 17278 6840 20038 6896
rect 17217 6838 20038 6840
rect 17217 6835 17283 6838
rect 19238 6808 20038 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 8477 6354 8543 6357
rect 8845 6354 8911 6357
rect 8477 6352 8911 6354
rect 8477 6296 8482 6352
rect 8538 6296 8850 6352
rect 8906 6296 8911 6352
rect 8477 6294 8911 6296
rect 8477 6291 8543 6294
rect 8845 6291 8911 6294
rect 11145 6354 11211 6357
rect 17217 6354 17283 6357
rect 11145 6352 17283 6354
rect 11145 6296 11150 6352
rect 11206 6296 17222 6352
rect 17278 6296 17283 6352
rect 11145 6294 17283 6296
rect 11145 6291 11211 6294
rect 17217 6291 17283 6294
rect 18505 6218 18571 6221
rect 19238 6218 20038 6248
rect 18505 6216 20038 6218
rect 18505 6160 18510 6216
rect 18566 6160 20038 6216
rect 18505 6158 20038 6160
rect 18505 6155 18571 6158
rect 19238 6128 20038 6158
rect 8017 6082 8083 6085
rect 8753 6082 8819 6085
rect 8017 6080 8819 6082
rect 8017 6024 8022 6080
rect 8078 6024 8758 6080
rect 8814 6024 8819 6080
rect 8017 6022 8819 6024
rect 8017 6019 8083 6022
rect 8753 6019 8819 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 10409 3090 10475 3093
rect 11145 3090 11211 3093
rect 10409 3088 11211 3090
rect 10409 3032 10414 3088
rect 10470 3032 11150 3088
rect 11206 3032 11211 3088
rect 10409 3030 11211 3032
rect 10409 3027 10475 3030
rect 11145 3027 11211 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 19072 4528 19632
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 19616 5188 19632
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _386_
timestamp -25199
transform -1 0 4324 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp -25199
transform -1 0 4968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _388_
timestamp -25199
transform -1 0 5244 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _389_
timestamp -25199
transform 1 0 3312 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _390_
timestamp -25199
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _391_
timestamp -25199
transform -1 0 2852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _392_
timestamp -25199
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _393_
timestamp -25199
transform 1 0 9292 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp -25199
transform 1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _395_
timestamp -25199
transform 1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _396_
timestamp -25199
transform 1 0 6440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp -25199
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _398_
timestamp -25199
transform -1 0 14352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _399_
timestamp -25199
transform 1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _400_
timestamp -25199
transform -1 0 17664 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _401_
timestamp -25199
transform -1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _402_
timestamp -25199
transform -1 0 17664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _403_
timestamp -25199
transform -1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _404_
timestamp -25199
transform -1 0 17940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _405_
timestamp -25199
transform -1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp -25199
transform -1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp -25199
transform -1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp -25199
transform -1 0 16100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _409_
timestamp -25199
transform 1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _410_
timestamp -25199
transform -1 0 13524 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _411_
timestamp -25199
transform -1 0 13800 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _412_
timestamp -25199
transform -1 0 12420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _413_
timestamp -25199
transform -1 0 13616 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp -25199
transform -1 0 13892 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp -25199
transform -1 0 2300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _416_
timestamp -25199
transform -1 0 3496 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _417_
timestamp -25199
transform -1 0 2852 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _418_
timestamp -25199
transform -1 0 2852 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _419_
timestamp -25199
transform -1 0 2208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _420_
timestamp -25199
transform 1 0 2484 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _421_
timestamp -25199
transform 1 0 1840 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _422_
timestamp -25199
transform -1 0 3128 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _423_
timestamp -25199
transform -1 0 3588 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _424_
timestamp -25199
transform 1 0 2300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _425_
timestamp -25199
transform 1 0 8648 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _426_
timestamp -25199
transform -1 0 8740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor4_4  _427_
timestamp -25199
transform -1 0 11224 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _428_
timestamp -25199
transform 1 0 11224 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _429_
timestamp -25199
transform -1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _430_
timestamp -25199
transform 1 0 17940 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _431_
timestamp -25199
transform -1 0 18308 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp -25199
transform 1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _433_
timestamp -25199
transform 1 0 17664 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _434_
timestamp -25199
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _435_
timestamp -25199
transform 1 0 17388 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _436_
timestamp -25199
transform 1 0 13708 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _437_
timestamp -25199
transform 1 0 17664 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _438_
timestamp -25199
transform 1 0 14444 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__or3_4  _439_
timestamp -25199
transform -1 0 16284 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_4  _440_
timestamp -25199
transform 1 0 14076 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__or4_4  _441_
timestamp -25199
transform -1 0 16468 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _442_
timestamp -25199
transform 1 0 14904 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _443_
timestamp -25199
transform 1 0 14168 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _444_
timestamp -25199
transform 1 0 14536 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _445_
timestamp -25199
transform 1 0 14996 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_1  _446_
timestamp -25199
transform 1 0 14076 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _447_
timestamp -25199
transform 1 0 14444 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _448_
timestamp -25199
transform 1 0 14352 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _449_
timestamp -25199
transform -1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _450_
timestamp -25199
transform 1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _451_
timestamp -25199
transform -1 0 15640 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _452_
timestamp -25199
transform 1 0 15364 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _453_
timestamp -25199
transform -1 0 15180 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _454_
timestamp -25199
transform -1 0 15364 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_4  _455_
timestamp -25199
transform 1 0 14904 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__and2_1  _456_
timestamp -25199
transform -1 0 16468 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _457_
timestamp -25199
transform 1 0 16652 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _458_
timestamp -25199
transform -1 0 16560 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _459_
timestamp -25199
transform -1 0 15732 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _460_
timestamp -25199
transform 1 0 15548 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _461_
timestamp -25199
transform 1 0 18124 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _462_
timestamp -25199
transform 1 0 17940 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _463_
timestamp -25199
transform -1 0 17664 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _464_
timestamp -25199
transform -1 0 16560 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _465_
timestamp -25199
transform 1 0 17204 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _466_
timestamp -25199
transform 1 0 16652 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _467_
timestamp -25199
transform -1 0 17940 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _468_
timestamp -25199
transform -1 0 18124 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _469_
timestamp -25199
transform -1 0 18032 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _470_
timestamp -25199
transform -1 0 17572 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _471_
timestamp -25199
transform 1 0 16652 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _472_
timestamp -25199
transform -1 0 16008 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _473_
timestamp -25199
transform -1 0 17940 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _474_
timestamp -25199
transform 1 0 17204 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _475_
timestamp -25199
transform -1 0 18124 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _476_
timestamp -25199
transform 1 0 16836 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _477_
timestamp -25199
transform -1 0 17020 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _478_
timestamp -25199
transform 1 0 16836 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _479_
timestamp -25199
transform 1 0 15916 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _480_
timestamp -25199
transform 1 0 15364 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _481_
timestamp -25199
transform -1 0 18124 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _482_
timestamp -25199
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _483_
timestamp -25199
transform -1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _484_
timestamp -25199
transform 1 0 16836 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _485_
timestamp -25199
transform 1 0 16744 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _486_
timestamp -25199
transform 1 0 15272 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _487_
timestamp -25199
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _488_
timestamp -25199
transform -1 0 18492 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_4  _489_
timestamp -25199
transform -1 0 17480 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _490_
timestamp -25199
transform -1 0 17020 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _491_
timestamp -25199
transform 1 0 16560 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _492_
timestamp -25199
transform -1 0 16376 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _493_
timestamp -25199
transform 1 0 15640 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _494_
timestamp -25199
transform -1 0 16652 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _495_
timestamp -25199
transform 1 0 16652 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _496_
timestamp -25199
transform -1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _497_
timestamp -25199
transform -1 0 17664 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _498_
timestamp -25199
transform 1 0 14996 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _499_
timestamp -25199
transform 1 0 15180 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _500_
timestamp -25199
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _501_
timestamp -25199
transform -1 0 10396 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _502_
timestamp -25199
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _503_
timestamp -25199
transform 1 0 8004 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _504_
timestamp -25199
transform 1 0 9660 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _505_
timestamp -25199
transform 1 0 7084 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _506_
timestamp -25199
transform -1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _507_
timestamp -25199
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _508_
timestamp -25199
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _509_
timestamp -25199
transform 1 0 7636 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _510_
timestamp -25199
transform 1 0 8648 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _511_
timestamp -25199
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _512_
timestamp -25199
transform 1 0 3128 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _513_
timestamp -25199
transform 1 0 2300 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _514_
timestamp -25199
transform 1 0 1932 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _515_
timestamp -25199
transform 1 0 3772 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _516_
timestamp -25199
transform 1 0 3220 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _517_
timestamp -25199
transform 1 0 1472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _518_
timestamp -25199
transform 1 0 2300 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _519_
timestamp -25199
transform 1 0 2208 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _520_
timestamp -25199
transform -1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _521_
timestamp -25199
transform 1 0 2576 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _522_
timestamp -25199
transform -1 0 3220 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _523_
timestamp -25199
transform -1 0 2668 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _524_
timestamp -25199
transform 1 0 1656 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _525_
timestamp -25199
transform -1 0 4692 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _526_
timestamp -25199
transform 1 0 4140 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _527_
timestamp -25199
transform -1 0 4140 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _528_
timestamp -25199
transform 1 0 2668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _529_
timestamp -25199
transform -1 0 2300 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _530_
timestamp -25199
transform 1 0 2300 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _531_
timestamp -25199
transform 1 0 3312 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _532_
timestamp -25199
transform 1 0 1840 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _533_
timestamp -25199
transform 1 0 3036 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _534_
timestamp -25199
transform -1 0 2668 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _535_
timestamp -25199
transform 1 0 2668 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _536_
timestamp -25199
transform 1 0 3220 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _537_
timestamp -25199
transform 1 0 3772 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _538_
timestamp -25199
transform 1 0 3772 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _539_
timestamp -25199
transform 1 0 4600 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _540_
timestamp -25199
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _541_
timestamp -25199
transform 1 0 3956 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _542_
timestamp -25199
transform -1 0 3588 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _543_
timestamp -25199
transform 1 0 3588 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21ba_1  _544_
timestamp -25199
transform -1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _545_
timestamp -25199
transform -1 0 5060 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _546_
timestamp -25199
transform -1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _547_
timestamp -25199
transform 1 0 16284 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _548_
timestamp -25199
transform -1 0 16284 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _549_
timestamp -25199
transform -1 0 15364 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _550_
timestamp -25199
transform 1 0 15088 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _551_
timestamp -25199
transform -1 0 17112 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _552_
timestamp -25199
transform -1 0 15824 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _553_
timestamp -25199
transform 1 0 16008 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _554_
timestamp -25199
transform 1 0 10304 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _555_
timestamp -25199
transform 1 0 9292 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _556_
timestamp -25199
transform -1 0 10948 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _557_
timestamp -25199
transform -1 0 10764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _558_
timestamp -25199
transform 1 0 10764 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _559_
timestamp -25199
transform -1 0 16560 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _560_
timestamp -25199
transform -1 0 15824 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__or4_4  _561_
timestamp -25199
transform -1 0 15548 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _562_
timestamp -25199
transform 1 0 15180 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _563_
timestamp -25199
transform -1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_4  _564_
timestamp -25199
transform 1 0 15180 0 1 14144
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_1  _565_
timestamp -25199
transform 1 0 4508 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _566_
timestamp -25199
transform 1 0 4692 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _567_
timestamp -25199
transform -1 0 5612 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _568_
timestamp -25199
transform 1 0 5244 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _569_
timestamp -25199
transform -1 0 6256 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _570_
timestamp -25199
transform 1 0 6256 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _571_
timestamp -25199
transform 1 0 5704 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _572_
timestamp -25199
transform 1 0 6348 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _573_
timestamp -25199
transform 1 0 6348 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _574_
timestamp -25199
transform -1 0 6348 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _575_
timestamp -25199
transform -1 0 6440 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _576_
timestamp -25199
transform 1 0 5796 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _577_
timestamp -25199
transform 1 0 5520 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _578_
timestamp -25199
transform -1 0 6256 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _579_
timestamp -25199
transform 1 0 5980 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _580_
timestamp -25199
transform 1 0 5428 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _581_
timestamp -25199
transform 1 0 6992 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _582_
timestamp -25199
transform 1 0 6348 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _583_
timestamp -25199
transform 1 0 5060 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _584_
timestamp -25199
transform -1 0 5980 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _585_
timestamp -25199
transform 1 0 5152 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _586_
timestamp -25199
transform 1 0 5060 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _587_
timestamp -25199
transform 1 0 6624 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _588_
timestamp -25199
transform 1 0 5796 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _589_
timestamp -25199
transform -1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _590_
timestamp -25199
transform -1 0 6256 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _591_
timestamp -25199
transform -1 0 5152 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _592_
timestamp -25199
transform 1 0 4876 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _593_
timestamp -25199
transform -1 0 5796 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _594_
timestamp -25199
transform -1 0 4784 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _595_
timestamp -25199
transform -1 0 5152 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _596_
timestamp -25199
transform -1 0 5060 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _597_
timestamp -25199
transform -1 0 5520 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _598_
timestamp -25199
transform -1 0 5152 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _599_
timestamp -25199
transform 1 0 5336 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _600_
timestamp -25199
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _601_
timestamp -25199
transform 1 0 6164 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _602_
timestamp -25199
transform 1 0 6808 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _603_
timestamp -25199
transform -1 0 6992 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _604_
timestamp -25199
transform 1 0 6624 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _605_
timestamp -25199
transform -1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _606_
timestamp -25199
transform -1 0 9384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _607_
timestamp -25199
transform 1 0 8372 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _608_
timestamp -25199
transform 1 0 10488 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _609_
timestamp -25199
transform 1 0 9660 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _610_
timestamp -25199
transform 1 0 10120 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _611_
timestamp -25199
transform -1 0 13156 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _612_
timestamp -25199
transform 1 0 13156 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _613_
timestamp -25199
transform 1 0 12052 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _614_
timestamp -25199
transform -1 0 12696 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _615_
timestamp -25199
transform 1 0 11500 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _616_
timestamp -25199
transform -1 0 12512 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _617_
timestamp -25199
transform -1 0 12880 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _618_
timestamp -25199
transform -1 0 12880 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _619_
timestamp -25199
transform 1 0 14076 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _620_
timestamp -25199
transform 1 0 11960 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _621_
timestamp -25199
transform -1 0 12420 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _622_
timestamp -25199
transform -1 0 12512 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _623_
timestamp -25199
transform 1 0 11500 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _624_
timestamp -25199
transform -1 0 12236 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _625_
timestamp -25199
transform -1 0 12052 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _626_
timestamp -25199
transform 1 0 10580 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _627_
timestamp -25199
transform -1 0 11316 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _628_
timestamp -25199
transform 1 0 10120 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _629_
timestamp -25199
transform 1 0 10396 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _630_
timestamp -25199
transform 1 0 10764 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _631_
timestamp -25199
transform 1 0 10212 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _632_
timestamp -25199
transform -1 0 10120 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _633_
timestamp -25199
transform 1 0 11408 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _634_
timestamp -25199
transform -1 0 11408 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _635_
timestamp -25199
transform 1 0 10396 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _636_
timestamp -25199
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _637_
timestamp -25199
transform -1 0 9660 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _638_
timestamp -25199
transform 1 0 8924 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _639_
timestamp -25199
transform -1 0 10580 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _640_
timestamp -25199
transform 1 0 9936 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _641_
timestamp -25199
transform 1 0 10304 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _642_
timestamp -25199
transform -1 0 11040 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _643_
timestamp -25199
transform -1 0 10396 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _644_
timestamp -25199
transform -1 0 13064 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _645_
timestamp -25199
transform 1 0 9016 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _646_
timestamp -25199
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _647_
timestamp -25199
transform -1 0 9936 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _648_
timestamp -25199
transform -1 0 10672 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _649_
timestamp -25199
transform 1 0 10580 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _650_
timestamp -25199
transform 1 0 9936 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _651_
timestamp -25199
transform 1 0 10120 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _652_
timestamp -25199
transform 1 0 10580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _653_
timestamp -25199
transform -1 0 11316 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _654_
timestamp -25199
transform 1 0 11316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _655_
timestamp -25199
transform -1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _656_
timestamp -25199
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _657_
timestamp -25199
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _658_
timestamp -25199
transform 1 0 11868 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _659_
timestamp -25199
transform -1 0 13432 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _660_
timestamp -25199
transform -1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _661_
timestamp -25199
transform 1 0 13248 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _662_
timestamp -25199
transform -1 0 13524 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _663_
timestamp -25199
transform 1 0 12328 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _664_
timestamp -25199
transform -1 0 13616 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _665_
timestamp -25199
transform -1 0 12512 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _666_
timestamp -25199
transform 1 0 13248 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _667_
timestamp -25199
transform 1 0 13156 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _668_
timestamp -25199
transform 1 0 13892 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _669_
timestamp -25199
transform -1 0 13156 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _670_
timestamp -25199
transform -1 0 13800 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _671_
timestamp -25199
transform 1 0 13800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _672_
timestamp -25199
transform 1 0 12604 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _673_
timestamp -25199
transform 1 0 12144 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _674_
timestamp -25199
transform -1 0 14260 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _675_
timestamp -25199
transform -1 0 15548 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _676_
timestamp -25199
transform 1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _677_
timestamp -25199
transform -1 0 13892 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _678_
timestamp -25199
transform -1 0 13984 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _679_
timestamp -25199
transform 1 0 14628 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _680_
timestamp -25199
transform -1 0 15732 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _681_
timestamp -25199
transform 1 0 13892 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _682_
timestamp -25199
transform 1 0 13708 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _683_
timestamp -25199
transform 1 0 13708 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _684_
timestamp -25199
transform 1 0 13156 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _685_
timestamp -25199
transform 1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _686_
timestamp -25199
transform -1 0 13708 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _687_
timestamp -25199
transform -1 0 13708 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _688_
timestamp -25199
transform 1 0 14168 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _689_
timestamp -25199
transform 1 0 14076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _690_
timestamp -25199
transform -1 0 13892 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _691_
timestamp -25199
transform -1 0 13156 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _692_
timestamp -25199
transform 1 0 4416 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _693_
timestamp -25199
transform 1 0 4692 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _694_
timestamp -25199
transform 1 0 3864 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _695_
timestamp -25199
transform 1 0 1656 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _696_
timestamp -25199
transform 1 0 2208 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _697_
timestamp -25199
transform 1 0 1472 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _698_
timestamp -25199
transform 1 0 2852 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _699_
timestamp -25199
transform 1 0 4416 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _700_
timestamp -25199
transform 1 0 4416 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _701_
timestamp -25199
transform -1 0 5336 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _702_
timestamp -25199
transform 1 0 2208 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _703_
timestamp -25199
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _704_
timestamp -25199
transform -1 0 4324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _705_
timestamp -25199
transform 1 0 4140 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _706_
timestamp -25199
transform 1 0 3864 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _707_
timestamp -25199
transform 1 0 5152 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _708_
timestamp -25199
transform 1 0 5428 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_1  _709_
timestamp -25199
transform 1 0 8004 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _710_
timestamp -25199
transform 1 0 10212 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _711_
timestamp -25199
transform -1 0 8004 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _712_
timestamp -25199
transform -1 0 7084 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _713_
timestamp -25199
transform 1 0 6716 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _714_
timestamp -25199
transform 1 0 6992 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _715_
timestamp -25199
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _716_
timestamp -25199
transform -1 0 10212 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _717_
timestamp -25199
transform -1 0 9936 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _718_
timestamp -25199
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _719_
timestamp -25199
transform -1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _720_
timestamp -25199
transform -1 0 9016 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _721_
timestamp -25199
transform 1 0 8004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _722_
timestamp -25199
transform 1 0 3956 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _723_
timestamp -25199
transform -1 0 8004 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _724_
timestamp -25199
transform 1 0 8280 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _725_
timestamp -25199
transform -1 0 8280 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _726_
timestamp -25199
transform 1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _727_
timestamp -25199
transform -1 0 9292 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _728_
timestamp -25199
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _729_
timestamp -25199
transform -1 0 9292 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _730_
timestamp -25199
transform 1 0 9660 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _731_
timestamp -25199
transform 1 0 12696 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _732_
timestamp -25199
transform 1 0 12512 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _733_
timestamp -25199
transform -1 0 13156 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _734_
timestamp -25199
transform -1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _735_
timestamp -25199
transform 1 0 4324 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _736_
timestamp -25199
transform -1 0 4784 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _737_
timestamp -25199
transform 1 0 4784 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _738_
timestamp -25199
transform -1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _739_
timestamp -25199
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _740_
timestamp -25199
transform -1 0 6256 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _741_
timestamp -25199
transform -1 0 6624 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _742_
timestamp -25199
transform -1 0 9016 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _743_
timestamp -25199
transform -1 0 7820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _744_
timestamp -25199
transform -1 0 7728 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _745_
timestamp -25199
transform -1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _746_
timestamp -25199
transform -1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _747_
timestamp -25199
transform -1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _748_
timestamp -25199
transform -1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _749_
timestamp -25199
transform -1 0 6900 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _750_
timestamp -25199
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _751_
timestamp -25199
transform -1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _752_
timestamp -25199
transform -1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _753_
timestamp -25199
transform -1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _754_
timestamp -25199
transform -1 0 11316 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _755_
timestamp -25199
transform -1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _756_
timestamp -25199
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _757_
timestamp -25199
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _758_
timestamp -25199
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _759_
timestamp -25199
transform 1 0 13156 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _760_
timestamp -25199
transform 1 0 12236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _761_
timestamp -25199
transform 1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _762_
timestamp -25199
transform -1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _763_
timestamp -25199
transform 1 0 11776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _764_
timestamp -25199
transform 1 0 9660 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _765_
timestamp -25199
transform 1 0 11684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _766_
timestamp -25199
transform -1 0 13340 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _767_
timestamp -25199
transform -1 0 9200 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _768_
timestamp -25199
transform -1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _769_
timestamp -25199
transform 1 0 9384 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _770_
timestamp -25199
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _771_
timestamp -25199
transform -1 0 11316 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _772_
timestamp -25199
transform -1 0 3220 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _773_
timestamp -25199
transform 1 0 4324 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _774_
timestamp -25199
transform 1 0 5060 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _775_
timestamp -25199
transform 1 0 6808 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _776_
timestamp -25199
transform -1 0 8280 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _777_
timestamp -25199
transform 1 0 6348 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _778_
timestamp -25199
transform 1 0 6624 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _779_
timestamp -25199
transform 1 0 6440 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _780_
timestamp -25199
transform 1 0 5796 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _781_
timestamp -25199
transform 1 0 6348 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _782_
timestamp -25199
transform 1 0 4784 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _783_
timestamp -25199
transform 1 0 4416 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _784_
timestamp -25199
transform 1 0 4140 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _785_
timestamp -25199
transform 1 0 6532 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _786_
timestamp -25199
transform 1 0 6716 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _787_
timestamp -25199
transform 1 0 8556 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _788_
timestamp -25199
transform 1 0 10120 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _789_
timestamp -25199
transform 1 0 12696 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _790_
timestamp -25199
transform 1 0 12880 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _791_
timestamp -25199
transform 1 0 12604 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _792_
timestamp -25199
transform 1 0 12144 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _793_
timestamp -25199
transform 1 0 11224 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _794_
timestamp -25199
transform 1 0 11500 0 -1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _795_
timestamp -25199
transform 1 0 9476 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _796_
timestamp -25199
transform 1 0 11500 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _797_
timestamp -25199
transform 1 0 8924 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _798_
timestamp -25199
transform 1 0 10856 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _799_
timestamp -25199
transform -1 0 12236 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _800_
timestamp -25199
transform -1 0 9936 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _801_
timestamp -25199
transform 1 0 10212 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _802_
timestamp -25199
transform -1 0 10856 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _803_
timestamp -25199
transform 1 0 11776 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _804_
timestamp -25199
transform 1 0 9936 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 8004 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp -25199
transform -1 0 8832 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp -25199
transform 1 0 9568 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp -25199
transform -1 0 8280 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp -25199
transform 1 0 9568 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__bufinv_16  clkload0
timestamp -25199
transform 1 0 7084 0 -1 7616
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp -25199
transform 1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  clkload2
timestamp -25199
transform 1 0 6440 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_2  clone11
timestamp -25199
transform -1 0 8924 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout35
timestamp -25199
transform -1 0 13708 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp -25199
transform 1 0 10304 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout37
timestamp -25199
transform -1 0 11408 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp -25199
transform 1 0 11592 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout40
timestamp -25199
transform -1 0 8740 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp -25199
transform 1 0 10396 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout42
timestamp -25199
transform -1 0 5980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout43
timestamp -25199
transform 1 0 9476 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp -25199
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67
timestamp -25199
transform 1 0 7268 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73
timestamp -25199
transform 1 0 7820 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp -25199
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp -25199
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91
timestamp -25199
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp -25199
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636943256
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp -25199
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp -25199
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp -25199
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636943256
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636943256
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp -25199
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636943256
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_181
timestamp -25199
transform 1 0 17756 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp -25199
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636943256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636943256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636943256
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636943256
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp -25199
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp -25199
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp -25199
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp -25199
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_116
timestamp -25199
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_147
timestamp 1636943256
transform 1 0 14628 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_159
timestamp -25199
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp -25199
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636943256
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181
timestamp -25199
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp -25199
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636943256
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636943256
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -25199
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636943256
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp -25199
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_46
timestamp -25199
transform 1 0 5336 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_54
timestamp -25199
transform 1 0 6072 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_67
timestamp 1636943256
transform 1 0 7268 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_119
timestamp -25199
transform 1 0 12052 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_136
timestamp -25199
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636943256
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636943256
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636943256
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636943256
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_189
timestamp -25199
transform 1 0 18492 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636943256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636943256
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_27
timestamp -25199
transform 1 0 3588 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp -25199
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp -25199
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp -25199
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_82
timestamp 1636943256
transform 1 0 8648 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_94
timestamp -25199
transform 1 0 9752 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp -25199
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -25199
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_148
timestamp 1636943256
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_160
timestamp -25199
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636943256
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_181
timestamp -25199
transform 1 0 17756 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp -25199
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636943256
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636943256
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -25199
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_29
timestamp -25199
transform 1 0 3772 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_54
timestamp -25199
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_64
timestamp 1636943256
transform 1 0 6992 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_76
timestamp -25199
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_92
timestamp 1636943256
transform 1 0 9568 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_104
timestamp 1636943256
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_116
timestamp -25199
transform 1 0 11776 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_120
timestamp -25199
transform 1 0 12144 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_124
timestamp -25199
transform 1 0 12512 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_132
timestamp -25199
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp -25199
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636943256
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636943256
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1636943256
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1636943256
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_189
timestamp -25199
transform 1 0 18492 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636943256
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636943256
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_27
timestamp -25199
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_35
timestamp -25199
transform 1 0 4324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_48
timestamp -25199
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636943256
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_69
timestamp -25199
transform 1 0 7452 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_89
timestamp -25199
transform 1 0 9292 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp -25199
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp -25199
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp -25199
transform 1 0 11500 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp -25199
transform 1 0 11868 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_148
timestamp -25199
transform 1 0 14720 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_152
timestamp -25199
transform 1 0 15088 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp -25199
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1636943256
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_181
timestamp -25199
transform 1 0 17756 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_189
timestamp -25199
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636943256
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636943256
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp -25199
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_44
timestamp 1636943256
transform 1 0 5152 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_56
timestamp -25199
transform 1 0 6256 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_64
timestamp -25199
transform 1 0 6992 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_70
timestamp -25199
transform 1 0 7544 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp -25199
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_85
timestamp -25199
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_98
timestamp -25199
transform 1 0 10120 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_110
timestamp -25199
transform 1 0 11224 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_137
timestamp -25199
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_175
timestamp 1636943256
transform 1 0 17204 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636943256
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636943256
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_27
timestamp -25199
transform 1 0 3588 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp -25199
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp -25199
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp -25199
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp -25199
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_141
timestamp -25199
transform 1 0 14076 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_149
timestamp -25199
transform 1 0 14812 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_169
timestamp -25199
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636943256
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636943256
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -25199
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp -25199
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp -25199
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_124
timestamp -25199
transform 1 0 12512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp -25199
transform 1 0 13064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_134
timestamp -25199
transform 1 0 13432 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1636943256
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1636943256
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_165
timestamp -25199
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_189
timestamp -25199
transform 1 0 18492 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636943256
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_15
timestamp -25199
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_20
timestamp 1636943256
transform 1 0 2944 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_32
timestamp -25199
transform 1 0 4048 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_40
timestamp -25199
transform 1 0 4784 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp -25199
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp -25199
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_124
timestamp -25199
transform 1 0 12512 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_132
timestamp -25199
transform 1 0 13248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp -25199
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_164
timestamp -25199
transform 1 0 16192 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp -25199
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_20
timestamp -25199
transform 1 0 2944 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp -25199
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_29
timestamp -25199
transform 1 0 3772 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_45
timestamp -25199
transform 1 0 5244 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_63
timestamp -25199
transform 1 0 6900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -25199
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_89
timestamp -25199
transform 1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_102
timestamp -25199
transform 1 0 10488 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_131
timestamp -25199
transform 1 0 13156 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp -25199
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp -25199
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp -25199
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_43
timestamp -25199
transform 1 0 5060 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_49
timestamp -25199
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp -25199
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_70
timestamp -25199
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp -25199
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp -25199
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp -25199
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_119
timestamp 1636943256
transform 1 0 12052 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp -25199
transform 1 0 13156 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_146
timestamp 1636943256
transform 1 0 14536 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp -25199
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp -25199
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp -25199
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_22
timestamp -25199
transform 1 0 3128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_36
timestamp -25199
transform 1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_56
timestamp -25199
transform 1 0 6256 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_64
timestamp -25199
transform 1 0 6992 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp -25199
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_91
timestamp -25199
transform 1 0 9476 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_99
timestamp -25199
transform 1 0 10212 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_109
timestamp -25199
transform 1 0 11132 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_120
timestamp 1636943256
transform 1 0 12144 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_132
timestamp -25199
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1636943256
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1636943256
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_165
timestamp -25199
transform 1 0 16284 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_169
timestamp -25199
transform 1 0 16652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp -25199
transform 1 0 17020 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp -25199
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp -25199
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_18
timestamp -25199
transform 1 0 2760 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_36
timestamp 1636943256
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_48
timestamp -25199
transform 1 0 5520 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1636943256
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1636943256
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1636943256
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_93
timestamp -25199
transform 1 0 9660 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_97
timestamp -25199
transform 1 0 10028 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -25199
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_143
timestamp -25199
transform 1 0 14260 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_149
timestamp -25199
transform 1 0 14812 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp -25199
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_169
timestamp -25199
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_177
timestamp -25199
transform 1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_6
timestamp -25199
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_19
timestamp -25199
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp -25199
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp -25199
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_40
timestamp -25199
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_65
timestamp -25199
transform 1 0 7084 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp -25199
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_88
timestamp -25199
transform 1 0 9200 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_114
timestamp 1636943256
transform 1 0 11592 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_126
timestamp -25199
transform 1 0 12696 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp -25199
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_170
timestamp -25199
transform 1 0 16744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_177
timestamp -25199
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_188
timestamp -25199
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_6
timestamp -25199
transform 1 0 1656 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_19
timestamp 1636943256
transform 1 0 2852 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_39
timestamp -25199
transform 1 0 4692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp -25199
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp -25199
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp -25199
transform 1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_98
timestamp -25199
transform 1 0 10120 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp -25199
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_113
timestamp -25199
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp -25199
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_144
timestamp -25199
transform 1 0 14352 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp -25199
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp -25199
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp -25199
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp -25199
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp -25199
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_41
timestamp -25199
transform 1 0 4876 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_75
timestamp -25199
transform 1 0 8004 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp -25199
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_99
timestamp -25199
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_117
timestamp 1636943256
transform 1 0 11868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp -25199
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1636943256
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_153
timestamp -25199
transform 1 0 15180 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_16_173
timestamp -25199
transform 1 0 17020 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_179
timestamp -25199
transform 1 0 17572 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_183
timestamp -25199
transform 1 0 17940 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_6
timestamp -25199
transform 1 0 1656 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_13
timestamp 1636943256
transform 1 0 2300 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_25
timestamp -25199
transform 1 0 3404 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_36
timestamp 1636943256
transform 1 0 4416 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_48
timestamp -25199
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp -25199
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_65
timestamp -25199
transform 1 0 7084 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_98
timestamp -25199
transform 1 0 10120 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp -25199
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_144
timestamp -25199
transform 1 0 14352 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_152
timestamp -25199
transform 1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp -25199
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp -25199
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1636943256
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_181
timestamp -25199
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp -25199
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_6
timestamp -25199
transform 1 0 1656 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_10
timestamp -25199
transform 1 0 2024 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_22
timestamp -25199
transform 1 0 3128 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp -25199
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_48
timestamp -25199
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp -25199
transform 1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp -25199
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636943256
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp -25199
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_119
timestamp 1636943256
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp -25199
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp -25199
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp -25199
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636943256
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_180
timestamp -25199
transform 1 0 17664 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_186
timestamp -25199
transform 1 0 18216 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp -25199
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_27
timestamp -25199
transform 1 0 3588 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp -25199
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_69
timestamp -25199
transform 1 0 7452 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_75
timestamp 1636943256
transform 1 0 8004 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_87
timestamp -25199
transform 1 0 9108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp -25199
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp -25199
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -25199
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_113
timestamp -25199
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_118
timestamp 1636943256
transform 1 0 11960 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_130
timestamp -25199
transform 1 0 13064 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_136
timestamp -25199
transform 1 0 13616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_159
timestamp -25199
transform 1 0 15732 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_176
timestamp -25199
transform 1 0 17296 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp -25199
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp -25199
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_12
timestamp -25199
transform 1 0 2208 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_19
timestamp -25199
transform 1 0 2852 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp -25199
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_37
timestamp -25199
transform 1 0 4508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_45
timestamp -25199
transform 1 0 5244 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp -25199
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1636943256
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1636943256
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_165
timestamp -25199
transform 1 0 16284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_180
timestamp -25199
transform 1 0 17664 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_186
timestamp -25199
transform 1 0 18216 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp -25199
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_9
timestamp -25199
transform 1 0 1932 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_13
timestamp 1636943256
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_25
timestamp 1636943256
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_37
timestamp 1636943256
transform 1 0 4508 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_49
timestamp -25199
transform 1 0 5612 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp -25199
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_72
timestamp 1636943256
transform 1 0 7728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_84
timestamp -25199
transform 1 0 8832 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_90
timestamp -25199
transform 1 0 9384 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp -25199
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp -25199
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_119
timestamp -25199
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_142
timestamp -25199
transform 1 0 14168 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp -25199
transform 1 0 14904 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp -25199
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_21_174
timestamp -25199
transform 1 0 17112 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_189
timestamp -25199
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_6
timestamp -25199
transform 1 0 1656 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_18
timestamp -25199
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp -25199
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_44
timestamp -25199
transform 1 0 5152 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_52
timestamp -25199
transform 1 0 5888 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_78
timestamp -25199
transform 1 0 8280 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp -25199
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp -25199
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121
timestamp -25199
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp -25199
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1636943256
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp -25199
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_80
timestamp -25199
transform 1 0 8464 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp -25199
transform 1 0 9200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp -25199
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_136
timestamp 1636943256
transform 1 0 13616 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_148
timestamp -25199
transform 1 0 14720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp -25199
transform 1 0 15088 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp -25199
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_189
timestamp -25199
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp -25199
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_11
timestamp 1636943256
transform 1 0 2116 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp -25199
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp -25199
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp -25199
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_46
timestamp -25199
transform 1 0 5336 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_57
timestamp -25199
transform 1 0 6348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_78
timestamp -25199
transform 1 0 8280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp -25199
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_96
timestamp -25199
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_119
timestamp -25199
transform 1 0 12052 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_123
timestamp -25199
transform 1 0 12420 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_131
timestamp -25199
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp -25199
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_141
timestamp -25199
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_149
timestamp -25199
transform 1 0 14812 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_160
timestamp -25199
transform 1 0 15824 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_164
timestamp -25199
transform 1 0 16192 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_168
timestamp -25199
transform 1 0 16560 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_174
timestamp -25199
transform 1 0 17112 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_185
timestamp -25199
transform 1 0 18124 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_189
timestamp -25199
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp -25199
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1636943256
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_33
timestamp -25199
transform 1 0 4140 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1636943256
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_64
timestamp -25199
transform 1 0 6992 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp -25199
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp -25199
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_116
timestamp -25199
transform 1 0 11776 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_124
timestamp -25199
transform 1 0 12512 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_135
timestamp -25199
transform 1 0 13524 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_143
timestamp -25199
transform 1 0 14260 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_153
timestamp -25199
transform 1 0 15180 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp -25199
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1636943256
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_181
timestamp -25199
transform 1 0 17756 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_189
timestamp -25199
transform 1 0 18492 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp -25199
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_19
timestamp -25199
transform 1 0 2852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp -25199
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_29
timestamp -25199
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_35
timestamp -25199
transform 1 0 4324 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_62
timestamp 1636943256
transform 1 0 6808 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_74
timestamp -25199
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp -25199
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1636943256
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp -25199
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_104
timestamp 1636943256
transform 1 0 10672 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_116
timestamp -25199
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp -25199
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_148
timestamp -25199
transform 1 0 14720 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_167
timestamp 1636943256
transform 1 0 16468 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_179
timestamp -25199
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_187
timestamp -25199
transform 1 0 18308 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_3
timestamp -25199
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_39
timestamp -25199
transform 1 0 4692 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_47
timestamp -25199
transform 1 0 5428 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_57
timestamp -25199
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_61
timestamp -25199
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_86
timestamp -25199
transform 1 0 9016 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_90
timestamp -25199
transform 1 0 9384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_97
timestamp -25199
transform 1 0 10028 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_106
timestamp -25199
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp -25199
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_121
timestamp -25199
transform 1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_134
timestamp -25199
transform 1 0 13432 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp -25199
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp -25199
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1636943256
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_181
timestamp -25199
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_189
timestamp -25199
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp -25199
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_11
timestamp -25199
transform 1 0 2116 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_19
timestamp -25199
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_23
timestamp -25199
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp -25199
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_29
timestamp -25199
transform 1 0 3772 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_35
timestamp -25199
transform 1 0 4324 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_49
timestamp -25199
transform 1 0 5612 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_55
timestamp -25199
transform 1 0 6164 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_63
timestamp 1636943256
transform 1 0 6900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_75
timestamp -25199
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp -25199
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_114
timestamp 1636943256
transform 1 0 11592 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_126
timestamp 1636943256
transform 1 0 12696 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp -25199
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_144
timestamp -25199
transform 1 0 14352 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_158
timestamp 1636943256
transform 1 0 15640 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_170
timestamp 1636943256
transform 1 0 16744 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_182
timestamp -25199
transform 1 0 17848 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_13
timestamp 1636943256
transform 1 0 2300 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_25
timestamp -25199
transform 1 0 3404 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_31
timestamp -25199
transform 1 0 3956 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp -25199
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_60
timestamp 1636943256
transform 1 0 6624 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_72
timestamp 1636943256
transform 1 0 7728 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_84
timestamp -25199
transform 1 0 8832 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_93
timestamp -25199
transform 1 0 9660 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_101
timestamp -25199
transform 1 0 10396 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp -25199
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_123
timestamp -25199
transform 1 0 12420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_130
timestamp -25199
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_138
timestamp -25199
transform 1 0 13800 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_144
timestamp -25199
transform 1 0 14352 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1636943256
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_181
timestamp -25199
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_189
timestamp -25199
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1636943256
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1636943256
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp -25199
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp -25199
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_42
timestamp -25199
transform 1 0 4968 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_64
timestamp 1636943256
transform 1 0 6992 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp -25199
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_85
timestamp -25199
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_93
timestamp -25199
transform 1 0 9660 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_170
timestamp 1636943256
transform 1 0 16744 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_182
timestamp -25199
transform 1 0 17848 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1636943256
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1636943256
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp -25199
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_29
timestamp 1636943256
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_41
timestamp -25199
transform 1 0 4876 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_76
timestamp -25199
transform 1 0 8096 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_31_85
timestamp 1636943256
transform 1 0 8924 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_97
timestamp -25199
transform 1 0 10028 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_105
timestamp -25199
transform 1 0 10764 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp -25199
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1636943256
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_125
timestamp -25199
transform 1 0 12604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_139
timestamp -25199
transform 1 0 13892 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_141
timestamp -25199
transform 1 0 14076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_172
timestamp 1636943256
transform 1 0 16928 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_184
timestamp -25199
transform 1 0 18032 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input1
timestamp -25199
transform 1 0 7268 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp -25199
transform 1 0 1380 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp -25199
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -25199
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -25199
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp -25199
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp -25199
transform 1 0 9752 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp -25199
transform -1 0 18584 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp -25199
transform -1 0 16560 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -25199
transform -1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp -25199
transform -1 0 18584 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input12
timestamp -25199
transform 1 0 1380 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input13
timestamp -25199
transform -1 0 18584 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -25199
transform -1 0 18584 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp -25199
transform -1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp -25199
transform -1 0 18584 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp -25199
transform -1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp -25199
transform -1 0 18584 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp -25199
transform -1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp -25199
transform 1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp -25199
transform 1 0 12972 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input22
timestamp -25199
transform -1 0 16928 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp -25199
transform 1 0 6348 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input24
timestamp -25199
transform 1 0 14076 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp -25199
transform -1 0 16560 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp -25199
transform 1 0 1380 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp -25199
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp -25199
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp -25199
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp -25199
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp -25199
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp -25199
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp -25199
transform 1 0 1380 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  max_cap39
timestamp -25199
transform -1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp -25199
transform 1 0 1380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_32
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_33
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_34
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_35
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_36
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_37
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_38
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_39
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_40
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_41
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_42
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_43
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_44
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_45
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_46
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_47
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_48
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_49
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_50
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_51
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_52
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_53
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_54
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_55
timestamp -25199
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp -25199
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_56
timestamp -25199
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp -25199
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_57
timestamp -25199
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp -25199
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_58
timestamp -25199
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp -25199
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_59
timestamp -25199
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp -25199
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_60
timestamp -25199
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp -25199
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_61
timestamp -25199
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp -25199
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_62
timestamp -25199
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp -25199
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_63
timestamp -25199
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp -25199
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1
timestamp -25199
transform -1 0 2576 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer2
timestamp -25199
transform -1 0 17848 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  rebuffer3
timestamp -25199
transform 1 0 9292 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer4
timestamp -25199
transform -1 0 15456 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  rebuffer5
timestamp -25199
transform -1 0 16744 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer19
timestamp -25199
transform -1 0 6624 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer20
timestamp -25199
transform -1 0 5980 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer21
timestamp -25199
transform -1 0 4784 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  rebuffer22
timestamp -25199
transform -1 0 8188 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp -25199
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp -25199
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_70
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_71
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_72
timestamp -25199
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_74
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_75
timestamp -25199
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_77
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_78
timestamp -25199
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_79
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_80
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_81
timestamp -25199
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_83
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_84
timestamp -25199
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_86
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_87
timestamp -25199
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_89
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_90
timestamp -25199
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_92
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_93
timestamp -25199
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_95
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_96
timestamp -25199
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_97
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_98
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_99
timestamp -25199
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_101
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_102
timestamp -25199
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_103
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_104
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_105
timestamp -25199
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_106
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_107
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_108
timestamp -25199
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_110
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_111
timestamp -25199
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_113
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_114
timestamp -25199
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_116
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_117
timestamp -25199
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_119
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_120
timestamp -25199
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_121
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_122
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_123
timestamp -25199
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_124
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_125
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_126
timestamp -25199
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_127
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_128
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_129
timestamp -25199
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_130
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_131
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_132
timestamp -25199
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_133
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_134
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_135
timestamp -25199
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_136
timestamp -25199
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_137
timestamp -25199
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_138
timestamp -25199
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_139
timestamp -25199
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_140
timestamp -25199
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_141
timestamp -25199
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_142
timestamp -25199
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_143
timestamp -25199
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_144
timestamp -25199
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_145
timestamp -25199
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_146
timestamp -25199
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_147
timestamp -25199
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_148
timestamp -25199
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_149
timestamp -25199
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_150
timestamp -25199
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_151
timestamp -25199
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_152
timestamp -25199
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_153
timestamp -25199
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp -25199
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_155
timestamp -25199
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_156
timestamp -25199
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_157
timestamp -25199
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_158
timestamp -25199
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp -25199
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_160
timestamp -25199
transform 1 0 3680 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_161
timestamp -25199
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_162
timestamp -25199
transform 1 0 8832 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_163
timestamp -25199
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_164
timestamp -25199
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_165
timestamp -25199
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 19632 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 19632 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 out
port 3 nsew signal output
flabel metal2 s 6458 21382 6514 22182 0 FreeSans 224 90 0 0 psc[0]
port 4 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 psc[10]
port 5 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 psc[11]
port 6 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 psc[12]
port 7 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 psc[13]
port 8 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 psc[14]
port 9 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 psc[15]
port 10 nsew signal input
flabel metal3 s 19238 6128 20038 6248 0 FreeSans 480 0 0 0 psc[16]
port 11 nsew signal input
flabel metal3 s 19238 7488 20038 7608 0 FreeSans 480 0 0 0 psc[17]
port 12 nsew signal input
flabel metal3 s 19238 6808 20038 6928 0 FreeSans 480 0 0 0 psc[18]
port 13 nsew signal input
flabel metal3 s 19238 8848 20038 8968 0 FreeSans 480 0 0 0 psc[19]
port 14 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 psc[1]
port 15 nsew signal input
flabel metal3 s 19238 8168 20038 8288 0 FreeSans 480 0 0 0 psc[20]
port 16 nsew signal input
flabel metal3 s 19238 10888 20038 11008 0 FreeSans 480 0 0 0 psc[21]
port 17 nsew signal input
flabel metal3 s 19238 10208 20038 10328 0 FreeSans 480 0 0 0 psc[22]
port 18 nsew signal input
flabel metal3 s 19238 9528 20038 9648 0 FreeSans 480 0 0 0 psc[23]
port 19 nsew signal input
flabel metal3 s 19238 12248 20038 12368 0 FreeSans 480 0 0 0 psc[24]
port 20 nsew signal input
flabel metal3 s 19238 12928 20038 13048 0 FreeSans 480 0 0 0 psc[25]
port 21 nsew signal input
flabel metal3 s 19238 14288 20038 14408 0 FreeSans 480 0 0 0 psc[26]
port 22 nsew signal input
flabel metal3 s 19238 13608 20038 13728 0 FreeSans 480 0 0 0 psc[27]
port 23 nsew signal input
flabel metal2 s 12898 21382 12954 22182 0 FreeSans 224 90 0 0 psc[28]
port 24 nsew signal input
flabel metal2 s 14830 21382 14886 22182 0 FreeSans 224 90 0 0 psc[29]
port 25 nsew signal input
flabel metal2 s 5814 21382 5870 22182 0 FreeSans 224 90 0 0 psc[2]
port 26 nsew signal input
flabel metal2 s 13542 21382 13598 22182 0 FreeSans 224 90 0 0 psc[30]
port 27 nsew signal input
flabel metal2 s 14186 21382 14242 22182 0 FreeSans 224 90 0 0 psc[31]
port 28 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 psc[3]
port 29 nsew signal input
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 psc[4]
port 30 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 psc[5]
port 31 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 psc[6]
port 32 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 psc[7]
port 33 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 psc[8]
port 34 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 psc[9]
port 35 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 rst
port 36 nsew signal input
rlabel metal1 9982 19584 9982 19584 0 VGND
rlabel metal1 9982 19040 9982 19040 0 VPWR
rlabel metal2 4646 18462 4646 18462 0 _000_
rlabel metal1 4692 5814 4692 5814 0 _001_
rlabel metal1 4508 4250 4508 4250 0 _002_
rlabel metal1 6808 3706 6808 3706 0 _003_
rlabel metal1 7176 2618 7176 2618 0 _004_
rlabel metal2 8878 3230 8878 3230 0 _005_
rlabel metal2 10442 3774 10442 3774 0 _006_
rlabel metal1 12834 2958 12834 2958 0 _007_
rlabel metal1 13018 4046 13018 4046 0 _008_
rlabel metal1 12742 5134 12742 5134 0 _009_
rlabel metal1 12466 6392 12466 6392 0 _010_
rlabel metal1 5244 17850 5244 17850 0 _011_
rlabel metal1 11362 7786 11362 7786 0 _012_
rlabel metal1 11730 9486 11730 9486 0 _013_
rlabel metal1 9650 10234 9650 10234 0 _014_
rlabel metal1 11408 11662 11408 11662 0 _015_
rlabel metal2 9246 13464 9246 13464 0 _016_
rlabel metal1 11040 12954 11040 12954 0 _017_
rlabel metal2 12466 14688 12466 14688 0 _018_
rlabel metal2 9522 15844 9522 15844 0 _019_
rlabel metal2 10534 15708 10534 15708 0 _020_
rlabel metal1 10534 17544 10534 17544 0 _021_
rlabel metal2 7130 17374 7130 17374 0 _022_
rlabel metal2 12098 18530 12098 18530 0 _023_
rlabel metal1 10534 18394 10534 18394 0 _024_
rlabel metal1 7452 15538 7452 15538 0 _025_
rlabel metal1 6440 14926 6440 14926 0 _026_
rlabel metal1 6946 13192 6946 13192 0 _027_
rlabel metal1 6946 12104 6946 12104 0 _028_
rlabel metal1 5934 11050 5934 11050 0 _029_
rlabel metal1 6440 9690 6440 9690 0 _030_
rlabel metal1 5283 6970 5283 6970 0 _031_
rlabel metal1 2990 11186 2990 11186 0 _032_
rlabel metal2 2162 11288 2162 11288 0 _033_
rlabel metal2 6118 18836 6118 18836 0 _034_
rlabel metal2 6486 18564 6486 18564 0 _035_
rlabel metal1 8609 17238 8609 17238 0 _036_
rlabel metal1 7597 15402 7597 15402 0 _037_
rlabel metal1 7636 14042 7636 14042 0 _038_
rlabel metal1 7912 12954 7912 12954 0 _039_
rlabel metal1 8195 12138 8195 12138 0 _040_
rlabel metal1 7597 11050 7597 11050 0 _041_
rlabel metal1 8418 10234 8418 10234 0 _042_
rlabel metal1 6539 6698 6539 6698 0 _043_
rlabel metal1 6217 6358 6217 6358 0 _044_
rlabel metal1 5382 3706 5382 3706 0 _045_
rlabel metal1 8510 4148 8510 4148 0 _046_
rlabel metal2 8050 2856 8050 2856 0 _047_
rlabel via2 11178 3043 11178 3043 0 _048_
rlabel metal1 11592 3094 11592 3094 0 _049_
rlabel metal1 13892 2618 13892 2618 0 _050_
rlabel metal2 13846 3944 13846 3944 0 _051_
rlabel metal2 13662 5032 13662 5032 0 _052_
rlabel metal2 13478 6494 13478 6494 0 _053_
rlabel metal1 12328 7514 12328 7514 0 _054_
rlabel metal1 12144 9146 12144 9146 0 _055_
rlabel metal1 11231 9962 11231 9962 0 _056_
rlabel metal1 12091 11798 12091 11798 0 _057_
rlabel metal2 9798 13090 9798 13090 0 _058_
rlabel metal2 11822 13090 11822 13090 0 _059_
rlabel metal2 12834 14552 12834 14552 0 _060_
rlabel metal2 9062 15640 9062 15640 0 _061_
rlabel metal2 11638 15674 11638 15674 0 _062_
rlabel metal2 9522 17816 9522 17816 0 _063_
rlabel metal1 13577 18666 13577 18666 0 _064_
rlabel metal2 11270 18904 11270 18904 0 _065_
rlabel metal1 4784 16014 4784 16014 0 _066_
rlabel metal2 4646 16830 4646 16830 0 _067_
rlabel metal1 5198 16150 5198 16150 0 _068_
rlabel metal1 3220 12750 3220 12750 0 _069_
rlabel metal1 2438 12240 2438 12240 0 _070_
rlabel metal1 2576 10642 2576 10642 0 _071_
rlabel metal1 6256 7854 6256 7854 0 _072_
rlabel metal1 9476 7854 9476 7854 0 _073_
rlabel metal2 9982 7378 9982 7378 0 _074_
rlabel metal1 7774 6256 7774 6256 0 _075_
rlabel metal1 7176 8398 7176 8398 0 _076_
rlabel metal1 6532 8398 6532 8398 0 _077_
rlabel metal2 14306 17034 14306 17034 0 _078_
rlabel metal1 15410 12614 15410 12614 0 _079_
rlabel metal1 17480 13294 17480 13294 0 _080_
rlabel metal1 17342 12750 17342 12750 0 _081_
rlabel metal1 14134 12886 14134 12886 0 _082_
rlabel metal1 17480 10574 17480 10574 0 _083_
rlabel metal2 17250 10778 17250 10778 0 _084_
rlabel metal2 17158 10506 17158 10506 0 _085_
rlabel metal1 15824 7854 15824 7854 0 _086_
rlabel metal1 15870 7310 15870 7310 0 _087_
rlabel metal1 16192 7786 16192 7786 0 _088_
rlabel metal2 10534 8092 10534 8092 0 _089_
rlabel metal2 13386 17612 13386 17612 0 _090_
rlabel metal1 13248 18326 13248 18326 0 _091_
rlabel metal1 11914 17646 11914 17646 0 _092_
rlabel metal1 13386 15130 13386 15130 0 _093_
rlabel metal1 13570 14314 13570 14314 0 _094_
rlabel metal2 3174 17204 3174 17204 0 _095_
rlabel metal1 2346 17306 2346 17306 0 _096_
rlabel metal2 2622 16218 2622 16218 0 _097_
rlabel metal1 2208 12750 2208 12750 0 _098_
rlabel metal2 2714 12517 2714 12517 0 _099_
rlabel metal1 2254 9452 2254 9452 0 _100_
rlabel metal2 2622 8364 2622 8364 0 _101_
rlabel metal1 2842 8330 2842 8330 0 _102_
rlabel metal1 3082 7922 3082 7922 0 _103_
rlabel metal2 9890 6834 9890 6834 0 _104_
rlabel metal1 8510 5610 8510 5610 0 _105_
rlabel metal2 11178 6460 11178 6460 0 _106_
rlabel metal1 17434 7820 17434 7820 0 _107_
rlabel metal1 18032 9146 18032 9146 0 _108_
rlabel metal2 17250 9316 17250 9316 0 _109_
rlabel metal1 15502 12682 15502 12682 0 _110_
rlabel metal1 16146 12716 16146 12716 0 _111_
rlabel metal1 17756 8602 17756 8602 0 _112_
rlabel metal2 15778 11526 15778 11526 0 _113_
rlabel metal1 16974 13362 16974 13362 0 _114_
rlabel metal1 14582 12682 14582 12682 0 _115_
rlabel metal1 18078 14586 18078 14586 0 _116_
rlabel metal2 14950 14348 14950 14348 0 _117_
rlabel metal1 15456 17646 15456 17646 0 _118_
rlabel metal1 15364 18258 15364 18258 0 _119_
rlabel metal2 15778 18428 15778 18428 0 _120_
rlabel metal2 14950 17170 14950 17170 0 _121_
rlabel metal1 14590 18394 14590 18394 0 _122_
rlabel metal1 14950 18156 14950 18156 0 _123_
rlabel metal1 15916 17170 15916 17170 0 _124_
rlabel metal1 15134 17204 15134 17204 0 _125_
rlabel metal1 14674 16082 14674 16082 0 _126_
rlabel metal2 14674 16694 14674 16694 0 _127_
rlabel metal1 15410 17170 15410 17170 0 _128_
rlabel metal1 15916 17102 15916 17102 0 _129_
rlabel metal1 15824 17034 15824 17034 0 _130_
rlabel metal2 15410 16524 15410 16524 0 _131_
rlabel metal1 15180 15946 15180 15946 0 _132_
rlabel metal1 15686 16558 15686 16558 0 _133_
rlabel metal2 16238 16252 16238 16252 0 _134_
rlabel metal1 15945 16082 15945 16082 0 _135_
rlabel metal1 16514 12818 16514 12818 0 _136_
rlabel metal1 16054 13906 16054 13906 0 _137_
rlabel metal2 15134 13515 15134 13515 0 _138_
rlabel metal2 17066 14110 17066 14110 0 _139_
rlabel metal2 18446 14518 18446 14518 0 _140_
rlabel metal2 17986 14688 17986 14688 0 _141_
rlabel metal1 16882 15470 16882 15470 0 _142_
rlabel metal1 17158 15674 17158 15674 0 _143_
rlabel metal2 17618 15232 17618 15232 0 _144_
rlabel metal2 16698 14722 16698 14722 0 _145_
rlabel metal1 16882 14960 16882 14960 0 _146_
rlabel metal1 15594 15504 15594 15504 0 _147_
rlabel metal1 17158 15028 17158 15028 0 _148_
rlabel metal1 17204 14586 17204 14586 0 _149_
rlabel metal2 16698 15606 16698 15606 0 _150_
rlabel metal2 15962 15164 15962 15164 0 _151_
rlabel metal2 17342 6970 17342 6970 0 _152_
rlabel metal1 17710 10030 17710 10030 0 _153_
rlabel metal1 16422 10710 16422 10710 0 _154_
rlabel metal2 16882 11254 16882 11254 0 _155_
rlabel metal1 16422 11220 16422 11220 0 _156_
rlabel metal2 16422 10438 16422 10438 0 _157_
rlabel metal1 15134 10676 15134 10676 0 _158_
rlabel metal1 15456 10642 15456 10642 0 _159_
rlabel metal1 16652 10506 16652 10506 0 _160_
rlabel metal1 15778 10574 15778 10574 0 _161_
rlabel metal2 16330 9792 16330 9792 0 _162_
rlabel metal2 16882 8772 16882 8772 0 _163_
rlabel metal2 15502 9350 15502 9350 0 _164_
rlabel metal1 15594 9486 15594 9486 0 _165_
rlabel via1 15336 10098 15336 10098 0 _166_
rlabel metal1 17158 5678 17158 5678 0 _167_
rlabel metal2 16698 7667 16698 7667 0 _168_
rlabel metal2 16790 6290 16790 6290 0 _169_
rlabel metal1 16652 5202 16652 5202 0 _170_
rlabel metal1 16422 5338 16422 5338 0 _171_
rlabel metal2 15778 5916 15778 5916 0 _172_
rlabel metal2 16790 7548 16790 7548 0 _173_
rlabel metal2 15410 6732 15410 6732 0 _174_
rlabel metal1 14950 5746 14950 5746 0 _175_
rlabel metal1 16146 6358 16146 6358 0 _176_
rlabel metal1 15456 5882 15456 5882 0 _177_
rlabel metal1 16054 5066 16054 5066 0 _178_
rlabel metal1 16192 6426 16192 6426 0 _179_
rlabel metal1 10994 6324 10994 6324 0 _180_
rlabel metal1 10672 5882 10672 5882 0 _181_
rlabel metal1 9246 5066 9246 5066 0 _182_
rlabel metal1 10626 5202 10626 5202 0 _183_
rlabel metal1 7682 5780 7682 5780 0 _184_
rlabel metal2 9062 5508 9062 5508 0 _185_
rlabel metal2 9338 6052 9338 6052 0 _186_
rlabel metal1 7866 5644 7866 5644 0 _187_
rlabel metal1 8602 5270 8602 5270 0 _188_
rlabel metal1 10350 5270 10350 5270 0 _189_
rlabel metal1 3128 7514 3128 7514 0 _190_
rlabel metal1 4370 7786 4370 7786 0 _191_
rlabel metal2 4186 8364 4186 8364 0 _192_
rlabel metal1 3266 8976 3266 8976 0 _193_
rlabel metal1 4554 8942 4554 8942 0 _194_
rlabel metal1 3864 9010 3864 9010 0 _195_
rlabel metal1 2530 9588 2530 9588 0 _196_
rlabel metal1 4002 9418 4002 9418 0 _197_
rlabel metal1 3542 10778 3542 10778 0 _198_
rlabel metal2 1886 16252 1886 16252 0 _199_
rlabel metal1 3358 15878 3358 15878 0 _200_
rlabel metal1 2162 17204 2162 17204 0 _201_
rlabel metal1 2806 17238 2806 17238 0 _202_
rlabel metal1 2714 17136 2714 17136 0 _203_
rlabel metal1 4968 17782 4968 17782 0 _204_
rlabel metal1 3634 17068 3634 17068 0 _205_
rlabel metal1 2926 17170 2926 17170 0 _206_
rlabel metal2 3358 15980 3358 15980 0 _207_
rlabel metal2 2622 13566 2622 13566 0 _208_
rlabel metal1 3496 13294 3496 13294 0 _209_
rlabel metal2 4094 13804 4094 13804 0 _210_
rlabel metal1 4186 12886 4186 12886 0 _211_
rlabel metal2 4002 12988 4002 12988 0 _212_
rlabel metal2 2530 12240 2530 12240 0 _213_
rlabel metal1 3266 12104 3266 12104 0 _214_
rlabel metal1 3726 12410 3726 12410 0 _215_
rlabel metal1 4600 12750 4600 12750 0 _216_
rlabel metal2 4186 10812 4186 10812 0 _217_
rlabel metal1 4692 7922 4692 7922 0 _218_
rlabel metal2 4002 8330 4002 8330 0 _219_
rlabel metal1 4600 8058 4600 8058 0 _220_
rlabel metal1 3588 9554 3588 9554 0 _221_
rlabel metal2 4738 8908 4738 8908 0 _222_
rlabel metal1 5060 8466 5060 8466 0 _223_
rlabel metal2 9154 5712 9154 5712 0 _224_
rlabel metal1 15594 5134 15594 5134 0 _225_
rlabel metal1 15870 9996 15870 9996 0 _226_
rlabel metal1 15824 9690 15824 9690 0 _227_
rlabel metal1 15410 10030 15410 10030 0 _228_
rlabel metal1 16100 14042 16100 14042 0 _229_
rlabel metal1 16146 14586 16146 14586 0 _230_
rlabel metal2 15502 15198 15502 15198 0 _231_
rlabel metal2 16422 14620 16422 14620 0 _232_
rlabel metal1 10672 5338 10672 5338 0 _233_
rlabel metal1 10718 5678 10718 5678 0 _234_
rlabel metal2 10534 5882 10534 5882 0 _235_
rlabel metal1 11178 5644 11178 5644 0 _236_
rlabel via1 15341 14790 15341 14790 0 _237_
rlabel metal1 15640 5814 15640 5814 0 _238_
rlabel metal1 15180 5882 15180 5882 0 _239_
rlabel metal1 15318 14994 15318 14994 0 _240_
rlabel metal2 15870 14586 15870 14586 0 _241_
rlabel metal2 16238 12308 16238 12308 0 _242_
rlabel metal2 12558 14756 12558 14756 0 _243_
rlabel metal1 5228 17578 5228 17578 0 _244_
rlabel metal1 6348 16558 6348 16558 0 _245_
rlabel metal2 6210 17578 6210 17578 0 _246_
rlabel metal1 6348 16082 6348 16082 0 _247_
rlabel metal1 6716 15878 6716 15878 0 _248_
rlabel metal1 6072 14790 6072 14790 0 _249_
rlabel metal2 6026 14824 6026 14824 0 _250_
rlabel metal2 5934 13056 5934 13056 0 _251_
rlabel metal2 6394 13600 6394 13600 0 _252_
rlabel metal1 5980 12614 5980 12614 0 _253_
rlabel metal1 6762 12648 6762 12648 0 _254_
rlabel metal1 5152 10030 5152 10030 0 _255_
rlabel metal2 5566 11050 5566 11050 0 _256_
rlabel metal2 6026 9622 6026 9622 0 _257_
rlabel metal1 6548 9622 6548 9622 0 _258_
rlabel metal1 5566 7514 5566 7514 0 _259_
rlabel metal1 5382 8976 5382 8976 0 _260_
rlabel metal1 4876 7378 4876 7378 0 _261_
rlabel metal1 5244 5814 5244 5814 0 _262_
rlabel metal2 4738 6103 4738 6103 0 _263_
rlabel metal2 4738 4590 4738 4590 0 _264_
rlabel metal1 5198 4114 5198 4114 0 _265_
rlabel metal1 6164 3434 6164 3434 0 _266_
rlabel metal2 6210 3774 6210 3774 0 _267_
rlabel metal1 7130 2346 7130 2346 0 _268_
rlabel metal1 6532 2550 6532 2550 0 _269_
rlabel metal1 9062 3706 9062 3706 0 _270_
rlabel metal1 8802 3434 8802 3434 0 _271_
rlabel metal2 10534 3638 10534 3638 0 _272_
rlabel metal1 12926 3536 12926 3536 0 _273_
rlabel metal1 12466 4080 12466 4080 0 _274_
rlabel metal1 13018 2822 13018 2822 0 _275_
rlabel metal1 12098 3706 12098 3706 0 _276_
rlabel metal1 12039 6630 12039 6630 0 _277_
rlabel metal2 12374 4284 12374 4284 0 _278_
rlabel metal1 12328 5610 12328 5610 0 _279_
rlabel metal1 12466 5032 12466 5032 0 _280_
rlabel metal2 12006 6120 12006 6120 0 _281_
rlabel metal2 11546 7412 11546 7412 0 _282_
rlabel metal1 10810 7854 10810 7854 0 _283_
rlabel metal1 11316 8058 11316 8058 0 _284_
rlabel metal1 10626 9384 10626 9384 0 _285_
rlabel metal1 10442 9690 10442 9690 0 _286_
rlabel metal1 11316 10778 11316 10778 0 _287_
rlabel metal1 9982 10438 9982 10438 0 _288_
rlabel metal2 11822 11560 11822 11560 0 _289_
rlabel metal1 10409 14042 10409 14042 0 _290_
rlabel metal2 8694 13600 8694 13600 0 _291_
rlabel metal1 9200 12954 9200 12954 0 _292_
rlabel metal1 10626 12410 10626 12410 0 _293_
rlabel metal2 10350 13260 10350 13260 0 _294_
rlabel metal1 12880 14994 12880 14994 0 _295_
rlabel metal1 12650 14824 12650 14824 0 _296_
rlabel metal1 9568 15606 9568 15606 0 _297_
rlabel metal1 9233 15334 9233 15334 0 _298_
rlabel metal1 10120 16422 10120 16422 0 _299_
rlabel metal1 10350 15912 10350 15912 0 _300_
rlabel metal2 10534 17578 10534 17578 0 _301_
rlabel metal2 10718 17782 10718 17782 0 _302_
rlabel metal1 11684 17850 11684 17850 0 _303_
rlabel metal1 10948 18122 10948 18122 0 _304_
rlabel metal1 12374 16694 12374 16694 0 _305_
rlabel metal1 12788 17034 12788 17034 0 _306_
rlabel metal2 13478 17102 13478 17102 0 _307_
rlabel metal1 12880 16626 12880 16626 0 _308_
rlabel metal1 12880 16218 12880 16218 0 _309_
rlabel metal1 13018 15402 13018 15402 0 _310_
rlabel metal1 12742 13974 12742 13974 0 _311_
rlabel metal1 12646 14042 12646 14042 0 _312_
rlabel metal1 13064 13498 13064 13498 0 _313_
rlabel metal1 13386 13770 13386 13770 0 _314_
rlabel metal1 13662 13974 13662 13974 0 _315_
rlabel metal2 12558 12852 12558 12852 0 _316_
rlabel metal1 13340 11662 13340 11662 0 _317_
rlabel metal1 13616 10574 13616 10574 0 _318_
rlabel metal2 13202 10948 13202 10948 0 _319_
rlabel metal2 13386 10676 13386 10676 0 _320_
rlabel metal1 13754 10438 13754 10438 0 _321_
rlabel metal1 14306 7990 14306 7990 0 _322_
rlabel metal1 15088 8058 15088 8058 0 _323_
rlabel metal1 13708 7718 13708 7718 0 _324_
rlabel metal2 13294 7582 13294 7582 0 _325_
rlabel metal1 14168 7242 14168 7242 0 _326_
rlabel metal1 14306 7412 14306 7412 0 _327_
rlabel metal1 13984 7514 13984 7514 0 _328_
rlabel metal1 14260 8602 14260 8602 0 _329_
rlabel metal1 13616 10778 13616 10778 0 _330_
rlabel metal1 14030 11322 14030 11322 0 _331_
rlabel metal2 13938 11356 13938 11356 0 _332_
rlabel metal1 12834 10132 12834 10132 0 _333_
rlabel metal1 13156 8602 13156 8602 0 _334_
rlabel metal2 14214 9044 14214 9044 0 _335_
rlabel metal1 13984 9962 13984 9962 0 _336_
rlabel metal1 13156 10030 13156 10030 0 _337_
rlabel metal1 12673 10234 12673 10234 0 _338_
rlabel metal1 5014 14314 5014 14314 0 _339_
rlabel metal1 4830 15334 4830 15334 0 _340_
rlabel metal1 4876 14382 4876 14382 0 _341_
rlabel metal1 2254 14790 2254 14790 0 _342_
rlabel metal1 4094 14416 4094 14416 0 _343_
rlabel metal2 2898 15266 2898 15266 0 _344_
rlabel metal2 4370 15300 4370 15300 0 _345_
rlabel metal1 4922 15504 4922 15504 0 _346_
rlabel metal2 4830 15674 4830 15674 0 _347_
rlabel metal2 4554 15198 4554 15198 0 _348_
rlabel metal1 4462 15028 4462 15028 0 _349_
rlabel metal2 4002 14739 4002 14739 0 _350_
rlabel metal1 4462 14586 4462 14586 0 _351_
rlabel metal1 4922 14858 4922 14858 0 _352_
rlabel metal1 4968 12138 4968 12138 0 _353_
rlabel metal1 6532 11866 6532 11866 0 _354_
rlabel metal1 7958 7888 7958 7888 0 _355_
rlabel metal2 10166 6970 10166 6970 0 _356_
rlabel metal2 9246 8058 9246 8058 0 _357_
rlabel metal2 8188 7854 8188 7854 0 _358_
rlabel metal1 7866 7514 7866 7514 0 _359_
rlabel metal1 8096 8534 8096 8534 0 _360_
rlabel via1 8418 7854 8418 7854 0 _361_
rlabel metal1 8464 9078 8464 9078 0 _362_
rlabel metal1 9154 8908 9154 8908 0 _363_
rlabel metal1 9384 8602 9384 8602 0 _364_
rlabel metal1 8050 8840 8050 8840 0 _365_
rlabel metal1 9062 8534 9062 8534 0 _366_
rlabel metal1 8261 8942 8261 8942 0 _367_
rlabel metal2 9154 11356 9154 11356 0 _368_
rlabel metal1 5888 11526 5888 11526 0 _369_
rlabel metal2 8970 11084 8970 11084 0 _370_
rlabel metal2 8510 8262 8510 8262 0 _371_
rlabel metal1 7774 8058 7774 8058 0 _372_
rlabel metal2 8970 8092 8970 8092 0 _373_
rlabel metal2 9338 8500 9338 8500 0 _374_
rlabel metal1 8924 9146 8924 9146 0 _375_
rlabel metal1 9660 10778 9660 10778 0 _376_
rlabel metal1 9568 11186 9568 11186 0 _377_
rlabel metal1 12880 13430 12880 13430 0 _378_
rlabel metal1 12926 15504 12926 15504 0 _379_
rlabel metal1 12742 15334 12742 15334 0 _380_
rlabel metal2 4646 13702 4646 13702 0 _381_
rlabel metal2 5106 14756 5106 14756 0 _382_
rlabel metal1 4830 14790 4830 14790 0 _383_
rlabel metal1 6992 15130 6992 15130 0 _384_
rlabel metal2 9338 11356 9338 11356 0 _385_
rlabel metal3 1717 18428 1717 18428 0 clk
rlabel metal1 8924 14314 8924 14314 0 clknet_0_clk
rlabel metal2 7130 8908 7130 8908 0 clknet_2_0__leaf_clk
rlabel metal1 12604 5202 12604 5202 0 clknet_2_1__leaf_clk
rlabel metal1 5106 18700 5106 18700 0 clknet_2_2__leaf_clk
rlabel metal1 10902 18802 10902 18802 0 clknet_2_3__leaf_clk
rlabel metal1 5612 17306 5612 17306 0 counter\[0\]
rlabel metal2 4554 6562 4554 6562 0 counter\[10\]
rlabel metal1 7038 7412 7038 7412 0 counter\[11\]
rlabel metal1 8740 5202 8740 5202 0 counter\[12\]
rlabel metal2 8970 5746 8970 5746 0 counter\[13\]
rlabel metal2 9430 6290 9430 6290 0 counter\[14\]
rlabel via1 10057 7854 10057 7854 0 counter\[15\]
rlabel metal2 14858 7616 14858 7616 0 counter\[16\]
rlabel metal1 12558 4046 12558 4046 0 counter\[17\]
rlabel metal1 12236 6970 12236 6970 0 counter\[18\]
rlabel metal1 12282 6698 12282 6698 0 counter\[19\]
rlabel metal2 5750 17986 5750 17986 0 counter\[1\]
rlabel metal1 14122 8364 14122 8364 0 counter\[20\]
rlabel metal2 15594 10132 15594 10132 0 counter\[21\]
rlabel metal1 16422 11118 16422 11118 0 counter\[22\]
rlabel metal1 15594 11696 15594 11696 0 counter\[23\]
rlabel metal1 13478 13260 13478 13260 0 counter\[24\]
rlabel metal1 16376 13974 16376 13974 0 counter\[25\]
rlabel metal1 13846 14314 13846 14314 0 counter\[26\]
rlabel metal2 13570 15470 13570 15470 0 counter\[27\]
rlabel metal2 14398 16286 14398 16286 0 counter\[28\]
rlabel via1 15042 17187 15042 17187 0 counter\[29\]
rlabel metal2 1794 15232 1794 15232 0 counter\[2\]
rlabel metal1 12972 16966 12972 16966 0 counter\[30\]
rlabel metal1 13018 18224 13018 18224 0 counter\[31\]
rlabel metal2 2254 14654 2254 14654 0 counter\[3\]
rlabel metal1 6118 15436 6118 15436 0 counter\[4\]
rlabel metal1 6302 13906 6302 13906 0 counter\[5\]
rlabel metal2 7222 12614 7222 12614 0 counter\[6\]
rlabel metal1 5888 10642 5888 10642 0 counter\[7\]
rlabel metal1 6348 10030 6348 10030 0 counter\[8\]
rlabel metal1 6118 8466 6118 8466 0 counter\[9\]
rlabel metal1 2599 16626 2599 16626 0 net1
rlabel metal1 17342 6970 17342 6970 0 net10
rlabel metal2 18446 7310 18446 7310 0 net11
rlabel metal1 2576 16762 2576 16762 0 net12
rlabel metal1 17112 8466 17112 8466 0 net13
rlabel metal2 18354 10812 18354 10812 0 net14
rlabel metal1 17986 11118 17986 11118 0 net15
rlabel metal2 18354 9860 18354 9860 0 net16
rlabel metal1 17986 12206 17986 12206 0 net17
rlabel metal2 18446 12988 18446 12988 0 net18
rlabel metal1 18032 13906 18032 13906 0 net19
rlabel metal1 5934 7854 5934 7854 0 net2
rlabel metal1 18676 13838 18676 13838 0 net20
rlabel metal1 13202 16116 13202 16116 0 net21
rlabel metal2 14214 18190 14214 18190 0 net22
rlabel metal1 5198 16592 5198 16592 0 net23
rlabel metal1 13892 18394 13892 18394 0 net24
rlabel metal1 15410 18666 15410 18666 0 net25
rlabel metal1 1794 16524 1794 16524 0 net26
rlabel metal1 1978 13328 1978 13328 0 net27
rlabel metal1 2070 12852 2070 12852 0 net28
rlabel metal1 1610 12750 1610 12750 0 net29
rlabel metal1 2668 8262 2668 8262 0 net3
rlabel metal1 1610 9962 1610 9962 0 net30
rlabel metal2 1610 11220 1610 11220 0 net31
rlabel metal1 1702 9044 1702 9044 0 net32
rlabel metal1 2231 18190 2231 18190 0 net33
rlabel metal2 1426 12308 1426 12308 0 net34
rlabel metal1 5750 9622 5750 9622 0 net35
rlabel metal1 12466 2992 12466 2992 0 net36
rlabel metal1 6762 12852 6762 12852 0 net37
rlabel metal2 12006 13770 12006 13770 0 net38
rlabel metal1 16882 12818 16882 12818 0 net39
rlabel metal1 8740 6290 8740 6290 0 net4
rlabel metal1 8694 2822 8694 2822 0 net40
rlabel metal2 12650 5882 12650 5882 0 net41
rlabel metal1 6210 19380 6210 19380 0 net42
rlabel metal1 13754 18768 13754 18768 0 net43
rlabel metal1 1656 9554 1656 9554 0 net44
rlabel metal1 17434 8466 17434 8466 0 net45
rlabel metal1 10166 6732 10166 6732 0 net46
rlabel metal1 14720 19346 14720 19346 0 net47
rlabel metal1 15962 18938 15962 18938 0 net48
rlabel metal1 8464 5542 8464 5542 0 net5
rlabel metal2 5842 17000 5842 17000 0 net54
rlabel metal1 10166 6256 10166 6256 0 net6
rlabel metal1 4186 9588 4186 9588 0 net62
rlabel metal1 5382 10030 5382 10030 0 net63
rlabel metal1 4416 9010 4416 9010 0 net64
rlabel metal2 7406 9452 7406 9452 0 net65
rlabel metal1 9936 2550 9936 2550 0 net7
rlabel metal1 17848 6290 17848 6290 0 net8
rlabel metal2 17158 7616 17158 7616 0 net9
rlabel metal3 751 12988 751 12988 0 out
rlabel metal1 6946 19346 6946 19346 0 psc[0]
rlabel metal3 1050 8228 1050 8228 0 psc[10]
rlabel metal3 751 7548 751 7548 0 psc[11]
rlabel metal2 7774 1554 7774 1554 0 psc[12]
rlabel metal2 8418 1588 8418 1588 0 psc[13]
rlabel metal2 9062 1554 9062 1554 0 psc[14]
rlabel metal2 9706 1588 9706 1588 0 psc[15]
rlabel via2 18538 6205 18538 6205 0 psc[16]
rlabel metal1 16514 7344 16514 7344 0 psc[17]
rlabel metal2 17250 6817 17250 6817 0 psc[18]
rlabel metal2 18446 8721 18446 8721 0 psc[19]
rlabel metal3 751 15708 751 15708 0 psc[1]
rlabel metal1 18584 5678 18584 5678 0 psc[20]
rlabel metal2 18538 11033 18538 11033 0 psc[21]
rlabel metal2 18262 10693 18262 10693 0 psc[22]
rlabel via2 18538 9571 18538 9571 0 psc[23]
rlabel metal2 18538 12257 18538 12257 0 psc[24]
rlabel metal2 18538 13141 18538 13141 0 psc[25]
rlabel via2 18262 14365 18262 14365 0 psc[26]
rlabel metal2 18538 14025 18538 14025 0 psc[27]
rlabel metal1 12972 19278 12972 19278 0 psc[28]
rlabel metal2 16882 20026 16882 20026 0 psc[29]
rlabel metal1 6118 19278 6118 19278 0 psc[2]
rlabel metal1 13984 18258 13984 18258 0 psc[30]
rlabel metal1 16514 19380 16514 19380 0 psc[31]
rlabel metal3 751 15028 751 15028 0 psc[3]
rlabel metal3 751 14348 751 14348 0 psc[4]
rlabel metal3 751 11628 751 11628 0 psc[5]
rlabel metal3 751 12308 751 12308 0 psc[6]
rlabel metal3 1050 9588 1050 9588 0 psc[7]
rlabel metal3 751 10268 751 10268 0 psc[8]
rlabel metal3 751 8908 751 8908 0 psc[9]
rlabel metal3 1050 17748 1050 17748 0 rst
<< properties >>
string FIXED_BBOX 0 0 20038 22182
<< end >>
