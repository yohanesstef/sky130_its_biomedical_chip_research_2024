magic
tech sky130A
magscale 1 2
timestamp 1730101407
<< checkpaint >>
rect -3932 -1804 14137 16281
<< viali >>
rect 3617 9537 3651 9571
rect 3985 9537 4019 9571
rect 5273 9537 5307 9571
rect 5641 9537 5675 9571
rect 6101 9537 6135 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 7021 9537 7055 9571
rect 5549 9469 5583 9503
rect 3525 9401 3559 9435
rect 5825 9401 5859 9435
rect 5917 9401 5951 9435
rect 3801 9333 3835 9367
rect 5365 9333 5399 9367
rect 5457 9333 5491 9367
rect 6745 9333 6779 9367
rect 6929 9333 6963 9367
rect 2237 9129 2271 9163
rect 5549 9129 5583 9163
rect 1593 9061 1627 9095
rect 3157 9061 3191 9095
rect 3525 9061 3559 9095
rect 7021 9061 7055 9095
rect 2145 8993 2179 9027
rect 2513 8993 2547 9027
rect 3249 8993 3283 9027
rect 3893 8993 3927 9027
rect 4721 8993 4755 9027
rect 1409 8925 1443 8959
rect 2053 8925 2087 8959
rect 2697 8925 2731 8959
rect 2789 8925 2823 8959
rect 3028 8925 3062 8959
rect 3985 8925 4019 8959
rect 4813 8925 4847 8959
rect 5365 8925 5399 8959
rect 5549 8925 5583 8959
rect 5917 8925 5951 8959
rect 6009 8925 6043 8959
rect 6469 8925 6503 8959
rect 6653 8925 6687 8959
rect 6745 8925 6779 8959
rect 7389 8925 7423 8959
rect 7757 8925 7791 8959
rect 2881 8857 2915 8891
rect 2421 8789 2455 8823
rect 2513 8789 2547 8823
rect 4353 8789 4387 8823
rect 5181 8789 5215 8823
rect 5733 8789 5767 8823
rect 6193 8789 6227 8823
rect 6561 8789 6595 8823
rect 7205 8789 7239 8823
rect 8401 8789 8435 8823
rect 2421 8585 2455 8619
rect 5089 8517 5123 8551
rect 5457 8517 5491 8551
rect 6561 8517 6595 8551
rect 1409 8449 1443 8483
rect 1869 8449 1903 8483
rect 1961 8449 1995 8483
rect 2145 8449 2179 8483
rect 2237 8449 2271 8483
rect 2513 8449 2547 8483
rect 2605 8449 2639 8483
rect 2789 8449 2823 8483
rect 3341 8449 3375 8483
rect 3434 8449 3468 8483
rect 3525 8449 3559 8483
rect 3643 8449 3677 8483
rect 3801 8449 3835 8483
rect 3893 8449 3927 8483
rect 4077 8449 4111 8483
rect 4261 8449 4295 8483
rect 4445 8449 4479 8483
rect 5273 8449 5307 8483
rect 5733 8449 5767 8483
rect 6377 8449 6411 8483
rect 6653 8449 6687 8483
rect 6745 8449 6779 8483
rect 7665 8449 7699 8483
rect 8217 8449 8251 8483
rect 4169 8381 4203 8415
rect 4629 8381 4663 8415
rect 7757 8381 7791 8415
rect 8033 8381 8067 8415
rect 2145 8313 2179 8347
rect 2237 8313 2271 8347
rect 3157 8313 3191 8347
rect 5641 8313 5675 8347
rect 7481 8313 7515 8347
rect 1593 8245 1627 8279
rect 2789 8245 2823 8279
rect 6929 8245 6963 8279
rect 2329 8041 2363 8075
rect 7757 8041 7791 8075
rect 8401 8041 8435 8075
rect 1685 7905 1719 7939
rect 2789 7905 2823 7939
rect 7389 7905 7423 7939
rect 1409 7837 1443 7871
rect 2513 7837 2547 7871
rect 2605 7837 2639 7871
rect 2697 7837 2731 7871
rect 3065 7837 3099 7871
rect 5549 7837 5583 7871
rect 6469 7837 6503 7871
rect 6837 7837 6871 7871
rect 7021 7837 7055 7871
rect 7205 7837 7239 7871
rect 7297 7837 7331 7871
rect 7573 7837 7607 7871
rect 7849 7837 7883 7871
rect 8217 7837 8251 7871
rect 6653 7769 6687 7803
rect 8033 7769 8067 7803
rect 8125 7769 8159 7803
rect 3157 7701 3191 7735
rect 5641 7701 5675 7735
rect 1869 7497 1903 7531
rect 2053 7497 2087 7531
rect 3617 7429 3651 7463
rect 1501 7361 1535 7395
rect 1655 7361 1689 7395
rect 1961 7361 1995 7395
rect 2789 7361 2823 7395
rect 2881 7361 2915 7395
rect 3157 7361 3191 7395
rect 3249 7361 3283 7395
rect 3397 7361 3431 7395
rect 3525 7361 3559 7395
rect 3714 7361 3748 7395
rect 4077 7361 4111 7395
rect 4261 7361 4295 7395
rect 4629 7361 4663 7395
rect 5365 7361 5399 7395
rect 5549 7361 5583 7395
rect 5917 7361 5951 7395
rect 6745 7361 6779 7395
rect 8401 7361 8435 7395
rect 2605 7293 2639 7327
rect 4353 7293 4387 7327
rect 4445 7293 4479 7327
rect 4813 7293 4847 7327
rect 5641 7293 5675 7327
rect 5733 7293 5767 7327
rect 8677 7293 8711 7327
rect 3893 7225 3927 7259
rect 3065 7157 3099 7191
rect 6101 7157 6135 7191
rect 6653 7157 6687 7191
rect 3157 6953 3191 6987
rect 7021 6885 7055 6919
rect 5825 6817 5859 6851
rect 7776 6817 7810 6851
rect 1777 6749 1811 6783
rect 1961 6749 1995 6783
rect 3065 6749 3099 6783
rect 5365 6749 5399 6783
rect 5457 6749 5491 6783
rect 5549 6749 5583 6783
rect 5733 6749 5767 6783
rect 6009 6749 6043 6783
rect 6377 6749 6411 6783
rect 6525 6749 6559 6783
rect 6745 6749 6779 6783
rect 6842 6749 6876 6783
rect 7573 6749 7607 6783
rect 8033 6749 8067 6783
rect 8125 6749 8159 6783
rect 8217 6749 8251 6783
rect 6193 6681 6227 6715
rect 6653 6681 6687 6715
rect 7113 6681 7147 6715
rect 7297 6681 7331 6715
rect 7849 6681 7883 6715
rect 1961 6613 1995 6647
rect 5181 6613 5215 6647
rect 7481 6613 7515 6647
rect 7665 6613 7699 6647
rect 8309 6613 8343 6647
rect 3617 6409 3651 6443
rect 3985 6409 4019 6443
rect 4077 6409 4111 6443
rect 4169 6409 4203 6443
rect 1593 6341 1627 6375
rect 1777 6341 1811 6375
rect 3801 6341 3835 6375
rect 7205 6341 7239 6375
rect 4629 6273 4663 6307
rect 4721 6273 4755 6307
rect 1869 6205 1903 6239
rect 2145 6205 2179 6239
rect 4813 6205 4847 6239
rect 4905 6205 4939 6239
rect 6929 6205 6963 6239
rect 4445 6137 4479 6171
rect 1409 6069 1443 6103
rect 4353 6069 4387 6103
rect 8677 6069 8711 6103
rect 2237 5865 2271 5899
rect 3157 5865 3191 5899
rect 3985 5865 4019 5899
rect 6009 5865 6043 5899
rect 8033 5865 8067 5899
rect 2421 5797 2455 5831
rect 7757 5797 7791 5831
rect 1869 5729 1903 5763
rect 4261 5729 4295 5763
rect 1777 5661 1811 5695
rect 3249 5661 3283 5695
rect 6285 5661 6319 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 7389 5661 7423 5695
rect 7481 5661 7515 5695
rect 7941 5661 7975 5695
rect 8585 5661 8619 5695
rect 2053 5593 2087 5627
rect 2253 5593 2287 5627
rect 3801 5593 3835 5627
rect 4017 5593 4051 5627
rect 4537 5593 4571 5627
rect 6193 5593 6227 5627
rect 1409 5525 1443 5559
rect 4169 5525 4203 5559
rect 6561 5525 6595 5559
rect 7205 5525 7239 5559
rect 5733 5321 5767 5355
rect 3617 5253 3651 5287
rect 4261 5253 4295 5287
rect 4445 5253 4479 5287
rect 6529 5253 6563 5287
rect 6745 5253 6779 5287
rect 7113 5253 7147 5287
rect 1501 5185 1535 5219
rect 1593 5185 1627 5219
rect 4353 5185 4387 5219
rect 1869 5117 1903 5151
rect 6837 5117 6871 5151
rect 1777 4981 1811 5015
rect 6377 4981 6411 5015
rect 6561 4981 6595 5015
rect 8585 4981 8619 5015
rect 3525 4777 3559 4811
rect 6009 4777 6043 4811
rect 6745 4777 6779 4811
rect 8217 4709 8251 4743
rect 2053 4641 2087 4675
rect 6561 4641 6595 4675
rect 1777 4573 1811 4607
rect 3985 4573 4019 4607
rect 5733 4573 5767 4607
rect 6469 4573 6503 4607
rect 6929 4573 6963 4607
rect 3893 4505 3927 4539
rect 5825 4505 5859 4539
rect 6041 4505 6075 4539
rect 5641 4437 5675 4471
rect 6193 4437 6227 4471
rect 5549 4233 5583 4267
rect 5841 4233 5875 4267
rect 3893 4165 3927 4199
rect 4109 4165 4143 4199
rect 4721 4165 4755 4199
rect 5181 4165 5215 4199
rect 5641 4165 5675 4199
rect 7021 4165 7055 4199
rect 7481 4165 7515 4199
rect 4353 4097 4387 4131
rect 4537 4097 4571 4131
rect 4813 4097 4847 4131
rect 4997 4097 5031 4131
rect 5089 4097 5123 4131
rect 5365 4097 5399 4131
rect 7665 4097 7699 4131
rect 7849 4097 7883 4131
rect 8209 4097 8243 4131
rect 8309 4097 8343 4131
rect 2329 4029 2363 4063
rect 2053 3961 2087 3995
rect 4905 3961 4939 3995
rect 1869 3893 1903 3927
rect 4077 3893 4111 3927
rect 4261 3893 4295 3927
rect 5825 3893 5859 3927
rect 6009 3893 6043 3927
rect 2034 3689 2068 3723
rect 3525 3689 3559 3723
rect 5917 3689 5951 3723
rect 8217 3689 8251 3723
rect 1777 3553 1811 3587
rect 4169 3553 4203 3587
rect 6745 3553 6779 3587
rect 3985 3485 4019 3519
rect 6285 3485 6319 3519
rect 6469 3485 6503 3519
rect 8309 3485 8343 3519
rect 3893 3417 3927 3451
rect 4445 3417 4479 3451
rect 6193 3417 6227 3451
rect 8401 3417 8435 3451
rect 4445 3145 4479 3179
rect 6469 3145 6503 3179
rect 5917 3077 5951 3111
rect 6193 3009 6227 3043
rect 6561 3009 6595 3043
rect 8677 3009 8711 3043
rect 8033 2805 8067 2839
rect 8309 2601 8343 2635
rect 8585 2397 8619 2431
<< metal1 >>
rect 1104 9818 9016 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 9016 9818
rect 1104 9744 9016 9766
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 5316 9676 5672 9704
rect 5316 9664 5322 9676
rect 3234 9596 3240 9648
rect 3292 9636 3298 9648
rect 3292 9608 4016 9636
rect 3292 9596 3298 9608
rect 3602 9528 3608 9580
rect 3660 9528 3666 9580
rect 3988 9577 4016 9608
rect 5644 9577 5672 9676
rect 3973 9571 4031 9577
rect 3973 9537 3985 9571
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 5629 9571 5687 9577
rect 5629 9537 5641 9571
rect 5675 9537 5687 9571
rect 5629 9531 5687 9537
rect 3418 9392 3424 9444
rect 3476 9432 3482 9444
rect 3513 9435 3571 9441
rect 3513 9432 3525 9435
rect 3476 9404 3525 9432
rect 3476 9392 3482 9404
rect 3513 9401 3525 9404
rect 3559 9432 3571 9435
rect 3970 9432 3976 9444
rect 3559 9404 3976 9432
rect 3559 9401 3571 9404
rect 3513 9395 3571 9401
rect 3970 9392 3976 9404
rect 4028 9392 4034 9444
rect 5276 9432 5304 9531
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 6089 9571 6147 9577
rect 6089 9568 6101 9571
rect 5868 9540 6101 9568
rect 5868 9528 5874 9540
rect 6089 9537 6101 9540
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6512 9540 6561 9568
rect 6512 9528 6518 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 7024 9500 7052 9531
rect 5592 9472 5948 9500
rect 5592 9460 5598 9472
rect 5626 9432 5632 9444
rect 5276 9404 5632 9432
rect 5626 9392 5632 9404
rect 5684 9432 5690 9444
rect 5920 9441 5948 9472
rect 6748 9472 7052 9500
rect 5813 9435 5871 9441
rect 5813 9432 5825 9435
rect 5684 9404 5825 9432
rect 5684 9392 5690 9404
rect 5813 9401 5825 9404
rect 5859 9401 5871 9435
rect 5813 9395 5871 9401
rect 5905 9435 5963 9441
rect 5905 9401 5917 9435
rect 5951 9401 5963 9435
rect 5905 9395 5963 9401
rect 3602 9324 3608 9376
rect 3660 9364 3666 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3660 9336 3801 9364
rect 3660 9324 3666 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 5350 9324 5356 9376
rect 5408 9324 5414 9376
rect 5445 9367 5503 9373
rect 5445 9333 5457 9367
rect 5491 9364 5503 9367
rect 5718 9364 5724 9376
rect 5491 9336 5724 9364
rect 5491 9333 5503 9336
rect 5445 9327 5503 9333
rect 5718 9324 5724 9336
rect 5776 9324 5782 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 6748 9373 6776 9472
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6696 9336 6745 9364
rect 6696 9324 6702 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 6917 9367 6975 9373
rect 6917 9333 6929 9367
rect 6963 9364 6975 9367
rect 7006 9364 7012 9376
rect 6963 9336 7012 9364
rect 6963 9333 6975 9336
rect 6917 9327 6975 9333
rect 7006 9324 7012 9336
rect 7064 9324 7070 9376
rect 1104 9274 9016 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 9016 9274
rect 1104 9200 9016 9222
rect 2222 9120 2228 9172
rect 2280 9120 2286 9172
rect 5537 9163 5595 9169
rect 2332 9132 2774 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 2332 9092 2360 9132
rect 1627 9064 2360 9092
rect 2746 9092 2774 9132
rect 5537 9129 5549 9163
rect 5583 9160 5595 9163
rect 5626 9160 5632 9172
rect 5583 9132 5632 9160
rect 5583 9129 5595 9132
rect 5537 9123 5595 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 3142 9092 3148 9104
rect 2746 9064 3148 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 2133 9027 2191 9033
rect 2133 8993 2145 9027
rect 2179 9024 2191 9027
rect 2332 9024 2360 9064
rect 3142 9052 3148 9064
rect 3200 9052 3206 9104
rect 3513 9095 3571 9101
rect 3513 9061 3525 9095
rect 3559 9092 3571 9095
rect 3559 9064 4752 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 2501 9027 2559 9033
rect 2501 9024 2513 9027
rect 2179 8996 2513 9024
rect 2179 8993 2191 8996
rect 2133 8987 2191 8993
rect 2501 8993 2513 8996
rect 2547 8993 2559 9027
rect 2501 8987 2559 8993
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 3237 9027 3295 9033
rect 2648 8996 2820 9024
rect 2648 8984 2654 8996
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 2792 8965 2820 8996
rect 3237 8993 3249 9027
rect 3283 9024 3295 9027
rect 3602 9024 3608 9036
rect 3283 8996 3608 9024
rect 3283 8993 3295 8996
rect 3237 8987 3295 8993
rect 3602 8984 3608 8996
rect 3660 8984 3666 9036
rect 4724 9033 4752 9064
rect 7006 9052 7012 9104
rect 7064 9052 7070 9104
rect 3881 9027 3939 9033
rect 3881 8993 3893 9027
rect 3927 8993 3939 9027
rect 3881 8987 3939 8993
rect 4709 9027 4767 9033
rect 4709 8993 4721 9027
rect 4755 9024 4767 9027
rect 4755 8996 5384 9024
rect 4755 8993 4767 8996
rect 4709 8987 4767 8993
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2087 8928 2697 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8956 2835 8959
rect 3016 8959 3074 8965
rect 3016 8956 3028 8959
rect 2823 8928 3028 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 3016 8925 3028 8928
rect 3062 8925 3074 8959
rect 3016 8919 3074 8925
rect 2700 8888 2728 8919
rect 2866 8888 2872 8900
rect 2424 8860 2636 8888
rect 2700 8860 2872 8888
rect 2424 8832 2452 8860
rect 2406 8780 2412 8832
rect 2464 8780 2470 8832
rect 2498 8780 2504 8832
rect 2556 8780 2562 8832
rect 2608 8820 2636 8860
rect 2866 8848 2872 8860
rect 2924 8848 2930 8900
rect 3234 8820 3240 8832
rect 2608 8792 3240 8820
rect 3234 8780 3240 8792
rect 3292 8820 3298 8832
rect 3896 8820 3924 8987
rect 5356 8968 5384 8996
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 6822 9024 6828 9036
rect 5776 8996 6040 9024
rect 5776 8984 5782 8996
rect 3970 8916 3976 8968
rect 4028 8916 4034 8968
rect 4798 8916 4804 8968
rect 4856 8916 4862 8968
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 6012 8965 6040 8996
rect 6472 8996 6828 9024
rect 6472 8965 6500 8996
rect 6822 8984 6828 8996
rect 6880 8984 6886 9036
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 5997 8959 6055 8965
rect 5997 8925 6009 8959
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8925 6515 8959
rect 6457 8919 6515 8925
rect 5920 8888 5948 8919
rect 6472 8888 6500 8919
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 6733 8959 6791 8965
rect 6733 8925 6745 8959
rect 6779 8956 6791 8959
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 6779 8928 7389 8956
rect 6779 8925 6791 8928
rect 6733 8919 6791 8925
rect 7377 8925 7389 8928
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 7745 8959 7803 8965
rect 7745 8925 7757 8959
rect 7791 8956 7803 8959
rect 8110 8956 8116 8968
rect 7791 8928 8116 8956
rect 7791 8925 7803 8928
rect 7745 8919 7803 8925
rect 5736 8860 6500 8888
rect 3292 8792 3924 8820
rect 3292 8780 3298 8792
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4341 8823 4399 8829
rect 4341 8820 4353 8823
rect 4304 8792 4353 8820
rect 4304 8780 4310 8792
rect 4341 8789 4353 8792
rect 4387 8789 4399 8823
rect 4341 8783 4399 8789
rect 5169 8823 5227 8829
rect 5169 8789 5181 8823
rect 5215 8820 5227 8823
rect 5442 8820 5448 8832
rect 5215 8792 5448 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 5736 8829 5764 8860
rect 5721 8823 5779 8829
rect 5721 8789 5733 8823
rect 5767 8789 5779 8823
rect 5721 8783 5779 8789
rect 6178 8780 6184 8832
rect 6236 8780 6242 8832
rect 6549 8823 6607 8829
rect 6549 8789 6561 8823
rect 6595 8820 6607 8823
rect 6748 8820 6776 8919
rect 8110 8916 8116 8928
rect 8168 8916 8174 8968
rect 6595 8792 6776 8820
rect 6595 8789 6607 8792
rect 6549 8783 6607 8789
rect 7190 8780 7196 8832
rect 7248 8780 7254 8832
rect 8202 8780 8208 8832
rect 8260 8820 8266 8832
rect 8389 8823 8447 8829
rect 8389 8820 8401 8823
rect 8260 8792 8401 8820
rect 8260 8780 8266 8792
rect 8389 8789 8401 8792
rect 8435 8789 8447 8823
rect 8389 8783 8447 8789
rect 1104 8730 9016 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 9016 8730
rect 1104 8656 9016 8678
rect 2406 8576 2412 8628
rect 2464 8576 2470 8628
rect 2498 8576 2504 8628
rect 2556 8616 2562 8628
rect 3326 8616 3332 8628
rect 2556 8588 3332 8616
rect 2556 8576 2562 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 4246 8616 4252 8628
rect 3717 8588 4252 8616
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1854 8440 1860 8492
rect 1912 8440 1918 8492
rect 1946 8440 1952 8492
rect 2004 8440 2010 8492
rect 2133 8483 2191 8489
rect 2133 8449 2145 8483
rect 2179 8449 2191 8483
rect 2133 8443 2191 8449
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2271 8452 2452 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2148 8412 2176 8443
rect 2148 8384 2268 8412
rect 2130 8304 2136 8356
rect 2188 8304 2194 8356
rect 2240 8353 2268 8384
rect 2225 8347 2283 8353
rect 2225 8313 2237 8347
rect 2271 8313 2283 8347
rect 2424 8344 2452 8452
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2590 8440 2596 8492
rect 2648 8440 2654 8492
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8480 2835 8483
rect 2958 8480 2964 8492
rect 2823 8452 2964 8480
rect 2823 8449 2835 8452
rect 2777 8443 2835 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3326 8440 3332 8492
rect 3384 8440 3390 8492
rect 3422 8483 3480 8489
rect 3422 8449 3434 8483
rect 3468 8449 3480 8483
rect 3422 8443 3480 8449
rect 3252 8412 3280 8440
rect 3437 8412 3465 8443
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 3631 8483 3689 8489
rect 3631 8449 3643 8483
rect 3677 8480 3689 8483
rect 3717 8480 3745 8588
rect 4246 8576 4252 8588
rect 4304 8576 4310 8628
rect 5460 8588 6776 8616
rect 5460 8560 5488 8588
rect 5077 8551 5135 8557
rect 5077 8548 5089 8551
rect 3896 8520 5089 8548
rect 3677 8452 3745 8480
rect 3677 8449 3689 8452
rect 3631 8443 3689 8449
rect 3786 8440 3792 8492
rect 3844 8440 3850 8492
rect 3896 8489 3924 8520
rect 5077 8517 5089 8520
rect 5123 8517 5135 8551
rect 5077 8511 5135 8517
rect 5442 8508 5448 8560
rect 5500 8508 5506 8560
rect 5552 8520 5856 8548
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 3252 8384 3465 8412
rect 4080 8356 4108 8443
rect 4246 8440 4252 8492
rect 4304 8440 4310 8492
rect 4338 8440 4344 8492
rect 4396 8480 4402 8492
rect 4433 8483 4491 8489
rect 4433 8480 4445 8483
rect 4396 8452 4445 8480
rect 4396 8440 4402 8452
rect 4433 8449 4445 8452
rect 4479 8480 4491 8483
rect 4522 8480 4528 8492
rect 4479 8452 4528 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5552 8480 5580 8520
rect 5307 8452 5580 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5626 8440 5632 8492
rect 5684 8480 5690 8492
rect 5721 8483 5779 8489
rect 5721 8480 5733 8483
rect 5684 8452 5733 8480
rect 5684 8440 5690 8452
rect 5721 8449 5733 8452
rect 5767 8449 5779 8483
rect 5828 8480 5856 8520
rect 6178 8508 6184 8560
rect 6236 8548 6242 8560
rect 6549 8551 6607 8557
rect 6549 8548 6561 8551
rect 6236 8520 6561 8548
rect 6236 8508 6242 8520
rect 6549 8517 6561 8520
rect 6595 8517 6607 8551
rect 6549 8511 6607 8517
rect 6270 8480 6276 8492
rect 5828 8452 6276 8480
rect 5721 8443 5779 8449
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4617 8415 4675 8421
rect 4617 8381 4629 8415
rect 4663 8412 4675 8415
rect 4663 8384 6316 8412
rect 4663 8381 4675 8384
rect 4617 8375 4675 8381
rect 3145 8347 3203 8353
rect 2424 8316 3096 8344
rect 2225 8307 2283 8313
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 1581 8279 1639 8285
rect 1581 8276 1593 8279
rect 1544 8248 1593 8276
rect 1544 8236 1550 8248
rect 1581 8245 1593 8248
rect 1627 8276 1639 8279
rect 2590 8276 2596 8288
rect 1627 8248 2596 8276
rect 1627 8245 1639 8248
rect 1581 8239 1639 8245
rect 2590 8236 2596 8248
rect 2648 8236 2654 8288
rect 2774 8236 2780 8288
rect 2832 8236 2838 8288
rect 3068 8276 3096 8316
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 3191 8316 3924 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 3510 8276 3516 8288
rect 3068 8248 3516 8276
rect 3510 8236 3516 8248
rect 3568 8236 3574 8288
rect 3896 8276 3924 8316
rect 4062 8304 4068 8356
rect 4120 8304 4126 8356
rect 4172 8276 4200 8375
rect 4798 8304 4804 8356
rect 4856 8344 4862 8356
rect 5442 8344 5448 8356
rect 4856 8316 5448 8344
rect 4856 8304 4862 8316
rect 5442 8304 5448 8316
rect 5500 8344 5506 8356
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5500 8316 5641 8344
rect 5500 8304 5506 8316
rect 5629 8313 5641 8316
rect 5675 8313 5687 8347
rect 5629 8307 5687 8313
rect 3896 8248 4200 8276
rect 6288 8276 6316 8384
rect 6380 8344 6408 8443
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6748 8489 6776 8588
rect 6641 8483 6699 8489
rect 6641 8480 6653 8483
rect 6512 8452 6653 8480
rect 6512 8440 6518 8452
rect 6641 8449 6653 8452
rect 6687 8449 6699 8483
rect 6641 8443 6699 8449
rect 6733 8483 6791 8489
rect 6733 8449 6745 8483
rect 6779 8449 6791 8483
rect 6733 8443 6791 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 7699 8452 8156 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 7742 8372 7748 8424
rect 7800 8372 7806 8424
rect 8018 8372 8024 8424
rect 8076 8372 8082 8424
rect 8128 8412 8156 8452
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 8386 8412 8392 8424
rect 8128 8384 8392 8412
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 6546 8344 6552 8356
rect 6380 8316 6552 8344
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 6656 8316 7420 8344
rect 6656 8276 6684 8316
rect 6288 8248 6684 8276
rect 6914 8236 6920 8288
rect 6972 8236 6978 8288
rect 7392 8276 7420 8316
rect 7466 8304 7472 8356
rect 7524 8304 7530 8356
rect 7558 8276 7564 8288
rect 7392 8248 7564 8276
rect 7558 8236 7564 8248
rect 7616 8236 7622 8288
rect 1104 8186 9016 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 9016 8186
rect 1104 8112 9016 8134
rect 1854 8032 1860 8084
rect 1912 8072 1918 8084
rect 2317 8075 2375 8081
rect 2317 8072 2329 8075
rect 1912 8044 2329 8072
rect 1912 8032 1918 8044
rect 2317 8041 2329 8044
rect 2363 8041 2375 8075
rect 2317 8035 2375 8041
rect 7742 8032 7748 8084
rect 7800 8032 7806 8084
rect 8386 8032 8392 8084
rect 8444 8032 8450 8084
rect 1673 7939 1731 7945
rect 1673 7905 1685 7939
rect 1719 7936 1731 7939
rect 1719 7908 2728 7936
rect 1719 7905 1731 7908
rect 1673 7899 1731 7905
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1854 7828 1860 7880
rect 1912 7868 1918 7880
rect 2501 7871 2559 7877
rect 2501 7868 2513 7871
rect 1912 7840 2513 7868
rect 1912 7828 1918 7840
rect 2501 7837 2513 7840
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2590 7828 2596 7880
rect 2648 7828 2654 7880
rect 2700 7877 2728 7908
rect 2774 7896 2780 7948
rect 2832 7896 2838 7948
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 7377 7939 7435 7945
rect 7377 7936 7389 7939
rect 6972 7908 7389 7936
rect 6972 7896 6978 7908
rect 7377 7905 7389 7908
rect 7423 7905 7435 7939
rect 7377 7899 7435 7905
rect 7484 7908 7880 7936
rect 2685 7871 2743 7877
rect 2685 7837 2697 7871
rect 2731 7868 2743 7871
rect 2958 7868 2964 7880
rect 2731 7840 2964 7868
rect 2731 7837 2743 7840
rect 2685 7831 2743 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3142 7868 3148 7880
rect 3099 7840 3148 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 5534 7828 5540 7880
rect 5592 7828 5598 7880
rect 6178 7828 6184 7880
rect 6236 7868 6242 7880
rect 6457 7871 6515 7877
rect 6457 7868 6469 7871
rect 6236 7840 6469 7868
rect 6236 7828 6242 7840
rect 6457 7837 6469 7840
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6871 7840 7021 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 7282 7828 7288 7880
rect 7340 7868 7346 7880
rect 7484 7868 7512 7908
rect 7340 7840 7512 7868
rect 7340 7828 7346 7840
rect 7558 7828 7564 7880
rect 7616 7828 7622 7880
rect 7852 7877 7880 7908
rect 8018 7896 8024 7948
rect 8076 7896 8082 7948
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 8036 7868 8064 7896
rect 8036 7840 8156 7868
rect 7837 7831 7895 7837
rect 6546 7760 6552 7812
rect 6604 7800 6610 7812
rect 6641 7803 6699 7809
rect 6641 7800 6653 7803
rect 6604 7772 6653 7800
rect 6604 7760 6610 7772
rect 6641 7769 6653 7772
rect 6687 7769 6699 7803
rect 7208 7800 7236 7828
rect 8128 7809 8156 7840
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 8021 7803 8079 7809
rect 8021 7800 8033 7803
rect 7208 7772 8033 7800
rect 6641 7763 6699 7769
rect 8021 7769 8033 7772
rect 8067 7769 8079 7803
rect 8021 7763 8079 7769
rect 8113 7803 8171 7809
rect 8113 7769 8125 7803
rect 8159 7800 8171 7803
rect 8570 7800 8576 7812
rect 8159 7772 8576 7800
rect 8159 7769 8171 7772
rect 8113 7763 8171 7769
rect 8570 7760 8576 7772
rect 8628 7760 8634 7812
rect 2866 7692 2872 7744
rect 2924 7732 2930 7744
rect 3145 7735 3203 7741
rect 3145 7732 3157 7735
rect 2924 7704 3157 7732
rect 2924 7692 2930 7704
rect 3145 7701 3157 7704
rect 3191 7701 3203 7735
rect 3145 7695 3203 7701
rect 5629 7735 5687 7741
rect 5629 7701 5641 7735
rect 5675 7732 5687 7735
rect 5902 7732 5908 7744
rect 5675 7704 5908 7732
rect 5675 7701 5687 7704
rect 5629 7695 5687 7701
rect 5902 7692 5908 7704
rect 5960 7692 5966 7744
rect 1104 7642 9016 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 9016 7642
rect 1104 7568 9016 7590
rect 1854 7488 1860 7540
rect 1912 7488 1918 7540
rect 2041 7531 2099 7537
rect 2041 7497 2053 7531
rect 2087 7528 2099 7531
rect 2590 7528 2596 7540
rect 2087 7500 2596 7528
rect 2087 7497 2099 7500
rect 2041 7491 2099 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 3476 7500 4660 7528
rect 3476 7488 3482 7500
rect 1762 7420 1768 7472
rect 1820 7460 1826 7472
rect 3605 7463 3663 7469
rect 3605 7460 3617 7463
rect 1820 7432 1992 7460
rect 1820 7420 1826 7432
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 1964 7401 1992 7432
rect 2884 7432 3617 7460
rect 2884 7404 2912 7432
rect 3605 7429 3617 7432
rect 3651 7429 3663 7463
rect 3605 7423 3663 7429
rect 1643 7395 1701 7401
rect 1643 7361 1655 7395
rect 1689 7392 1701 7395
rect 1949 7395 2007 7401
rect 1689 7364 1900 7392
rect 1689 7361 1701 7364
rect 1643 7355 1701 7361
rect 1872 7256 1900 7364
rect 1949 7361 1961 7395
rect 1995 7392 2007 7395
rect 2682 7392 2688 7404
rect 1995 7364 2688 7392
rect 1995 7361 2007 7364
rect 1949 7355 2007 7361
rect 2682 7352 2688 7364
rect 2740 7392 2746 7404
rect 2777 7395 2835 7401
rect 2777 7392 2789 7395
rect 2740 7364 2789 7392
rect 2740 7352 2746 7364
rect 2777 7361 2789 7364
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3418 7401 3424 7404
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7361 3295 7395
rect 3237 7355 3295 7361
rect 3385 7395 3424 7401
rect 3385 7361 3397 7395
rect 3385 7355 3424 7361
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 3252 7324 3280 7355
rect 3418 7352 3424 7355
rect 3476 7352 3482 7404
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 3702 7395 3760 7401
rect 3702 7392 3714 7395
rect 3620 7364 3714 7392
rect 3620 7336 3648 7364
rect 3702 7361 3714 7364
rect 3748 7361 3760 7395
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 3702 7355 3760 7361
rect 3896 7364 4077 7392
rect 2639 7296 3280 7324
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 3602 7284 3608 7336
rect 3660 7284 3666 7336
rect 3896 7265 3924 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4249 7395 4307 7401
rect 4249 7361 4261 7395
rect 4295 7392 4307 7395
rect 4522 7392 4528 7404
rect 4295 7364 4528 7392
rect 4295 7361 4307 7364
rect 4249 7355 4307 7361
rect 4522 7352 4528 7364
rect 4580 7352 4586 7404
rect 4632 7401 4660 7500
rect 5810 7460 5816 7472
rect 5368 7432 5816 7460
rect 5368 7401 5396 7432
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 5353 7395 5411 7401
rect 5353 7361 5365 7395
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7361 5595 7395
rect 5537 7355 5595 7361
rect 4341 7327 4399 7333
rect 4341 7293 4353 7327
rect 4387 7293 4399 7327
rect 4341 7287 4399 7293
rect 3881 7259 3939 7265
rect 1872 7228 2774 7256
rect 2746 7200 2774 7228
rect 3881 7225 3893 7259
rect 3927 7225 3939 7259
rect 4356 7256 4384 7287
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 5552 7324 5580 7355
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6638 7352 6644 7404
rect 6696 7392 6702 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6696 7364 6745 7392
rect 6696 7352 6702 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 8168 7364 8401 7392
rect 8168 7352 8174 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 4847 7296 5580 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 5626 7284 5632 7336
rect 5684 7284 5690 7336
rect 5721 7327 5779 7333
rect 5721 7293 5733 7327
rect 5767 7324 5779 7327
rect 6270 7324 6276 7336
rect 5767 7296 6276 7324
rect 5767 7293 5779 7296
rect 5721 7287 5779 7293
rect 5442 7256 5448 7268
rect 4356 7228 5448 7256
rect 3881 7219 3939 7225
rect 5442 7216 5448 7228
rect 5500 7216 5506 7268
rect 5534 7216 5540 7268
rect 5592 7256 5598 7268
rect 5736 7256 5764 7287
rect 6270 7284 6276 7296
rect 6328 7284 6334 7336
rect 8662 7284 8668 7336
rect 8720 7284 8726 7336
rect 5592 7228 5764 7256
rect 5592 7216 5598 7228
rect 2746 7160 2780 7200
rect 2774 7148 2780 7160
rect 2832 7188 2838 7200
rect 3053 7191 3111 7197
rect 3053 7188 3065 7191
rect 2832 7160 3065 7188
rect 2832 7148 2838 7160
rect 3053 7157 3065 7160
rect 3099 7157 3111 7191
rect 3053 7151 3111 7157
rect 3510 7148 3516 7200
rect 3568 7188 3574 7200
rect 4062 7188 4068 7200
rect 3568 7160 4068 7188
rect 3568 7148 3574 7160
rect 4062 7148 4068 7160
rect 4120 7188 4126 7200
rect 4430 7188 4436 7200
rect 4120 7160 4436 7188
rect 4120 7148 4126 7160
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 6089 7191 6147 7197
rect 6089 7157 6101 7191
rect 6135 7188 6147 7191
rect 6362 7188 6368 7200
rect 6135 7160 6368 7188
rect 6135 7157 6147 7160
rect 6089 7151 6147 7157
rect 6362 7148 6368 7160
rect 6420 7148 6426 7200
rect 6641 7191 6699 7197
rect 6641 7157 6653 7191
rect 6687 7188 6699 7191
rect 6730 7188 6736 7200
rect 6687 7160 6736 7188
rect 6687 7157 6699 7160
rect 6641 7151 6699 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 1104 7098 9016 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 9016 7098
rect 1104 7024 9016 7046
rect 3142 6944 3148 6996
rect 3200 6944 3206 6996
rect 2682 6876 2688 6928
rect 2740 6916 2746 6928
rect 3602 6916 3608 6928
rect 2740 6888 3608 6916
rect 2740 6876 2746 6888
rect 3602 6876 3608 6888
rect 3660 6876 3666 6928
rect 6178 6876 6184 6928
rect 6236 6916 6242 6928
rect 6546 6916 6552 6928
rect 6236 6888 6552 6916
rect 6236 6876 6242 6888
rect 6546 6876 6552 6888
rect 6604 6916 6610 6928
rect 7009 6919 7067 6925
rect 6604 6888 6868 6916
rect 6604 6876 6610 6888
rect 5810 6808 5816 6860
rect 5868 6808 5874 6860
rect 6012 6820 6776 6848
rect 1762 6740 1768 6792
rect 1820 6740 1826 6792
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 1964 6712 1992 6743
rect 2958 6740 2964 6792
rect 3016 6780 3022 6792
rect 3053 6783 3111 6789
rect 3053 6780 3065 6783
rect 3016 6752 3065 6780
rect 3016 6740 3022 6752
rect 3053 6749 3065 6752
rect 3099 6749 3111 6783
rect 3053 6743 3111 6749
rect 5258 6740 5264 6792
rect 5316 6780 5322 6792
rect 5353 6783 5411 6789
rect 5353 6780 5365 6783
rect 5316 6752 5365 6780
rect 5316 6740 5322 6752
rect 5353 6749 5365 6752
rect 5399 6749 5411 6783
rect 5353 6743 5411 6749
rect 5442 6740 5448 6792
rect 5500 6740 5506 6792
rect 5534 6740 5540 6792
rect 5592 6740 5598 6792
rect 5721 6783 5779 6789
rect 5721 6749 5733 6783
rect 5767 6780 5779 6783
rect 5902 6780 5908 6792
rect 5767 6752 5908 6780
rect 5767 6749 5779 6752
rect 5721 6743 5779 6749
rect 5902 6740 5908 6752
rect 5960 6740 5966 6792
rect 6012 6789 6040 6820
rect 6748 6792 6776 6820
rect 5997 6783 6055 6789
rect 5997 6749 6009 6783
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 6513 6783 6571 6789
rect 6513 6749 6525 6783
rect 6559 6780 6571 6783
rect 6559 6749 6592 6780
rect 6513 6743 6592 6749
rect 2774 6712 2780 6724
rect 1964 6684 2780 6712
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 6178 6672 6184 6724
rect 6236 6672 6242 6724
rect 1946 6604 1952 6656
rect 2004 6604 2010 6656
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5626 6644 5632 6656
rect 5215 6616 5632 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 6564 6644 6592 6743
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 6840 6789 6868 6888
rect 7009 6885 7021 6919
rect 7055 6885 7067 6919
rect 7009 6879 7067 6885
rect 6830 6783 6888 6789
rect 6830 6749 6842 6783
rect 6876 6749 6888 6783
rect 7024 6780 7052 6879
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 7764 6851 7822 6857
rect 7764 6848 7776 6851
rect 7248 6820 7776 6848
rect 7248 6808 7254 6820
rect 7764 6817 7776 6820
rect 7810 6817 7822 6851
rect 7764 6811 7822 6817
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7024 6752 7573 6780
rect 6830 6743 6888 6749
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7561 6743 7619 6749
rect 7668 6752 8033 6780
rect 6641 6715 6699 6721
rect 6641 6681 6653 6715
rect 6687 6712 6699 6715
rect 7098 6712 7104 6724
rect 6687 6684 7104 6712
rect 6687 6681 6699 6684
rect 6641 6675 6699 6681
rect 7098 6672 7104 6684
rect 7156 6672 7162 6724
rect 7285 6715 7343 6721
rect 7285 6681 7297 6715
rect 7331 6712 7343 6715
rect 7668 6712 7696 6752
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8021 6743 8079 6749
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8202 6740 8208 6792
rect 8260 6740 8266 6792
rect 7331 6684 7696 6712
rect 7331 6681 7343 6684
rect 7285 6675 7343 6681
rect 7300 6644 7328 6675
rect 7834 6672 7840 6724
rect 7892 6672 7898 6724
rect 6564 6616 7328 6644
rect 7469 6647 7527 6653
rect 7469 6613 7481 6647
rect 7515 6644 7527 6647
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 7515 6616 7665 6644
rect 7515 6613 7527 6616
rect 7469 6607 7527 6613
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 7653 6607 7711 6613
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 1104 6554 9016 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 9016 6554
rect 1104 6480 9016 6502
rect 2774 6440 2780 6452
rect 1596 6412 2780 6440
rect 1596 6381 1624 6412
rect 2774 6400 2780 6412
rect 2832 6440 2838 6452
rect 2832 6412 3464 6440
rect 2832 6400 2838 6412
rect 1581 6375 1639 6381
rect 1581 6341 1593 6375
rect 1627 6341 1639 6375
rect 1581 6335 1639 6341
rect 1762 6332 1768 6384
rect 1820 6332 1826 6384
rect 3142 6332 3148 6384
rect 3200 6332 3206 6384
rect 3436 6372 3464 6412
rect 3602 6400 3608 6452
rect 3660 6440 3666 6452
rect 3973 6443 4031 6449
rect 3973 6440 3985 6443
rect 3660 6412 3985 6440
rect 3660 6400 3666 6412
rect 3973 6409 3985 6412
rect 4019 6409 4031 6443
rect 3973 6403 4031 6409
rect 3789 6375 3847 6381
rect 3789 6372 3801 6375
rect 3436 6344 3801 6372
rect 3789 6341 3801 6344
rect 3835 6341 3847 6375
rect 3988 6372 4016 6403
rect 4062 6400 4068 6452
rect 4120 6400 4126 6452
rect 4157 6443 4215 6449
rect 4157 6409 4169 6443
rect 4203 6440 4215 6443
rect 4614 6440 4620 6452
rect 4203 6412 4620 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4614 6400 4620 6412
rect 4672 6440 4678 6452
rect 4890 6440 4896 6452
rect 4672 6412 4896 6440
rect 4672 6400 4678 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 3988 6344 4752 6372
rect 3789 6335 3847 6341
rect 1857 6239 1915 6245
rect 1857 6236 1869 6239
rect 1780 6208 1869 6236
rect 1780 6180 1808 6208
rect 1857 6205 1869 6208
rect 1903 6205 1915 6239
rect 1857 6199 1915 6205
rect 2130 6196 2136 6248
rect 2188 6196 2194 6248
rect 3804 6236 3832 6335
rect 4062 6264 4068 6316
rect 4120 6304 4126 6316
rect 4724 6313 4752 6344
rect 7190 6332 7196 6384
rect 7248 6332 7254 6384
rect 4617 6307 4675 6313
rect 4617 6304 4629 6307
rect 4120 6276 4629 6304
rect 4120 6264 4126 6276
rect 4617 6273 4629 6276
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 4801 6239 4859 6245
rect 3804 6208 4568 6236
rect 1762 6128 1768 6180
rect 1820 6128 1826 6180
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 4433 6171 4491 6177
rect 4433 6168 4445 6171
rect 4120 6140 4445 6168
rect 4120 6128 4126 6140
rect 4433 6137 4445 6140
rect 4479 6137 4491 6171
rect 4540 6168 4568 6208
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 4816 6168 4844 6199
rect 4890 6196 4896 6248
rect 4948 6196 4954 6248
rect 6914 6196 6920 6248
rect 6972 6196 6978 6248
rect 4540 6140 4844 6168
rect 4433 6131 4491 6137
rect 1397 6103 1455 6109
rect 1397 6069 1409 6103
rect 1443 6100 1455 6103
rect 2222 6100 2228 6112
rect 1443 6072 2228 6100
rect 1443 6069 1455 6072
rect 1397 6063 1455 6069
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 4341 6103 4399 6109
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 4706 6100 4712 6112
rect 4387 6072 4712 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 7926 6060 7932 6112
rect 7984 6100 7990 6112
rect 8665 6103 8723 6109
rect 8665 6100 8677 6103
rect 7984 6072 8677 6100
rect 7984 6060 7990 6072
rect 8665 6069 8677 6072
rect 8711 6069 8723 6103
rect 8665 6063 8723 6069
rect 1104 6010 9016 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 9016 6010
rect 1104 5936 9016 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 2225 5899 2283 5905
rect 2225 5896 2237 5899
rect 1544 5868 2237 5896
rect 1544 5856 1550 5868
rect 2225 5865 2237 5868
rect 2271 5896 2283 5899
rect 2271 5868 2774 5896
rect 2271 5865 2283 5868
rect 2225 5859 2283 5865
rect 2130 5788 2136 5840
rect 2188 5828 2194 5840
rect 2409 5831 2467 5837
rect 2409 5828 2421 5831
rect 2188 5800 2421 5828
rect 2188 5788 2194 5800
rect 2409 5797 2421 5800
rect 2455 5797 2467 5831
rect 2409 5791 2467 5797
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 1946 5760 1952 5772
rect 1903 5732 1952 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 1397 5559 1455 5565
rect 1397 5525 1409 5559
rect 1443 5556 1455 5559
rect 1578 5556 1584 5568
rect 1443 5528 1584 5556
rect 1443 5525 1455 5528
rect 1397 5519 1455 5525
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 1780 5556 1808 5655
rect 1964 5624 1992 5720
rect 2041 5627 2099 5633
rect 2041 5624 2053 5627
rect 1964 5596 2053 5624
rect 2041 5593 2053 5596
rect 2087 5593 2099 5627
rect 2041 5587 2099 5593
rect 2222 5584 2228 5636
rect 2280 5633 2286 5636
rect 2280 5627 2299 5633
rect 2287 5593 2299 5627
rect 2746 5624 2774 5868
rect 3142 5856 3148 5908
rect 3200 5856 3206 5908
rect 3973 5899 4031 5905
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4246 5896 4252 5908
rect 4019 5868 4252 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 5258 5896 5264 5908
rect 4948 5868 5264 5896
rect 4948 5856 4954 5868
rect 5258 5856 5264 5868
rect 5316 5896 5322 5908
rect 5997 5899 6055 5905
rect 5997 5896 6009 5899
rect 5316 5868 6009 5896
rect 5316 5856 5322 5868
rect 5997 5865 6009 5868
rect 6043 5865 6055 5899
rect 5997 5859 6055 5865
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7892 5868 8033 5896
rect 7892 5856 7898 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 7745 5831 7803 5837
rect 7745 5797 7757 5831
rect 7791 5828 7803 5831
rect 8294 5828 8300 5840
rect 7791 5800 8300 5828
rect 7791 5797 7803 5800
rect 7745 5791 7803 5797
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 4249 5763 4307 5769
rect 4249 5729 4261 5763
rect 4295 5760 4307 5763
rect 4614 5760 4620 5772
rect 4295 5732 4620 5760
rect 4295 5729 4307 5732
rect 4249 5723 4307 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 7006 5760 7012 5772
rect 6288 5732 7012 5760
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3694 5692 3700 5704
rect 3283 5664 3700 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 6288 5701 6316 5732
rect 7006 5720 7012 5732
rect 7064 5760 7070 5772
rect 8202 5760 8208 5772
rect 7064 5732 8208 5760
rect 7064 5720 7070 5732
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5661 6331 5695
rect 6273 5655 6331 5661
rect 6362 5652 6368 5704
rect 6420 5652 6426 5704
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 3789 5627 3847 5633
rect 3789 5624 3801 5627
rect 2746 5596 3801 5624
rect 2280 5587 2299 5593
rect 3789 5593 3801 5596
rect 3835 5624 3847 5627
rect 3878 5624 3884 5636
rect 3835 5596 3884 5624
rect 3835 5593 3847 5596
rect 3789 5587 3847 5593
rect 2280 5584 2286 5587
rect 3878 5584 3884 5596
rect 3936 5584 3942 5636
rect 4062 5633 4068 5636
rect 4005 5627 4068 5633
rect 4005 5593 4017 5627
rect 4051 5593 4068 5627
rect 4005 5587 4068 5593
rect 4062 5584 4068 5587
rect 4120 5584 4126 5636
rect 4525 5627 4583 5633
rect 4525 5624 4537 5627
rect 4172 5596 4537 5624
rect 3510 5556 3516 5568
rect 1780 5528 3516 5556
rect 3510 5516 3516 5528
rect 3568 5516 3574 5568
rect 4172 5565 4200 5596
rect 4525 5593 4537 5596
rect 4571 5593 4583 5627
rect 6181 5627 6239 5633
rect 6181 5624 6193 5627
rect 5750 5596 6193 5624
rect 4525 5587 4583 5593
rect 6181 5593 6193 5596
rect 6227 5593 6239 5627
rect 6564 5624 6592 5655
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 7466 5652 7472 5704
rect 7524 5652 7530 5704
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 7098 5624 7104 5636
rect 6564 5596 7104 5624
rect 6181 5587 6239 5593
rect 7098 5584 7104 5596
rect 7156 5624 7162 5636
rect 7742 5624 7748 5636
rect 7156 5596 7748 5624
rect 7156 5584 7162 5596
rect 7742 5584 7748 5596
rect 7800 5584 7806 5636
rect 4157 5559 4215 5565
rect 4157 5525 4169 5559
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 6546 5516 6552 5568
rect 6604 5516 6610 5568
rect 7190 5516 7196 5568
rect 7248 5516 7254 5568
rect 1104 5466 9016 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 9016 5466
rect 1104 5392 9016 5414
rect 5721 5355 5779 5361
rect 5721 5352 5733 5355
rect 3620 5324 5733 5352
rect 3620 5293 3648 5324
rect 5721 5321 5733 5324
rect 5767 5352 5779 5355
rect 6914 5352 6920 5364
rect 5767 5324 6920 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 6914 5312 6920 5324
rect 6972 5312 6978 5364
rect 3605 5287 3663 5293
rect 3605 5253 3617 5287
rect 3651 5253 3663 5287
rect 3605 5247 3663 5253
rect 4246 5244 4252 5296
rect 4304 5244 4310 5296
rect 4430 5244 4436 5296
rect 4488 5244 4494 5296
rect 6517 5287 6575 5293
rect 6517 5284 6529 5287
rect 4724 5256 6529 5284
rect 4724 5228 4752 5256
rect 6517 5253 6529 5256
rect 6563 5253 6575 5287
rect 6517 5247 6575 5253
rect 6733 5287 6791 5293
rect 6733 5253 6745 5287
rect 6779 5253 6791 5287
rect 6733 5247 6791 5253
rect 7101 5287 7159 5293
rect 7101 5253 7113 5287
rect 7147 5284 7159 5287
rect 7190 5284 7196 5296
rect 7147 5256 7196 5284
rect 7147 5253 7159 5256
rect 7101 5247 7159 5253
rect 1486 5176 1492 5228
rect 1544 5176 1550 5228
rect 1578 5176 1584 5228
rect 1636 5176 1642 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4706 5216 4712 5228
rect 4387 5188 4712 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 6178 5216 6184 5228
rect 5592 5188 6184 5216
rect 5592 5176 5598 5188
rect 6178 5176 6184 5188
rect 6236 5216 6242 5228
rect 6748 5216 6776 5247
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 6236 5188 6776 5216
rect 6236 5176 6242 5188
rect 1762 5108 1768 5160
rect 1820 5148 1826 5160
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1820 5120 1869 5148
rect 1820 5108 1826 5120
rect 1857 5117 1869 5120
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 5810 5108 5816 5160
rect 5868 5148 5874 5160
rect 5868 5120 6684 5148
rect 5868 5108 5874 5120
rect 6270 5040 6276 5092
rect 6328 5080 6334 5092
rect 6656 5080 6684 5120
rect 6822 5108 6828 5160
rect 6880 5108 6886 5160
rect 7466 5148 7472 5160
rect 6932 5120 7472 5148
rect 6932 5080 6960 5120
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 8220 5148 8248 5202
rect 8294 5148 8300 5160
rect 8220 5120 8300 5148
rect 8294 5108 8300 5120
rect 8352 5108 8358 5160
rect 6328 5052 6592 5080
rect 6656 5052 6960 5080
rect 6328 5040 6334 5052
rect 1765 5015 1823 5021
rect 1765 4981 1777 5015
rect 1811 5012 1823 5015
rect 2038 5012 2044 5024
rect 1811 4984 2044 5012
rect 1811 4981 1823 4984
rect 1765 4975 1823 4981
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 6564 5021 6592 5052
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 4981 6607 5015
rect 6549 4975 6607 4981
rect 8570 4972 8576 5024
rect 8628 4972 8634 5024
rect 1104 4922 9016 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 9016 4922
rect 1104 4848 9016 4870
rect 3510 4768 3516 4820
rect 3568 4768 3574 4820
rect 5997 4811 6055 4817
rect 5997 4777 6009 4811
rect 6043 4808 6055 4811
rect 6546 4808 6552 4820
rect 6043 4780 6552 4808
rect 6043 4777 6055 4780
rect 5997 4771 6055 4777
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 6733 4811 6791 4817
rect 6733 4777 6745 4811
rect 6779 4808 6791 4811
rect 7374 4808 7380 4820
rect 6779 4780 7380 4808
rect 6779 4777 6791 4780
rect 6733 4771 6791 4777
rect 7374 4768 7380 4780
rect 7432 4768 7438 4820
rect 6822 4700 6828 4752
rect 6880 4740 6886 4752
rect 8205 4743 8263 4749
rect 8205 4740 8217 4743
rect 6880 4712 8217 4740
rect 6880 4700 6886 4712
rect 8205 4709 8217 4712
rect 8251 4709 8263 4743
rect 8205 4703 8263 4709
rect 2038 4632 2044 4684
rect 2096 4632 2102 4684
rect 6546 4632 6552 4684
rect 6604 4632 6610 4684
rect 8570 4672 8576 4684
rect 6840 4644 8576 4672
rect 1762 4564 1768 4616
rect 1820 4564 1826 4616
rect 3694 4564 3700 4616
rect 3752 4604 3758 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3752 4576 3985 4604
rect 3752 4564 3758 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4604 5779 4607
rect 6362 4604 6368 4616
rect 5767 4576 6368 4604
rect 5767 4573 5779 4576
rect 5721 4567 5779 4573
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4604 6515 4607
rect 6840 4604 6868 4644
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 6503 4576 6868 4604
rect 6503 4573 6515 4576
rect 6457 4567 6515 4573
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 3881 4539 3939 4545
rect 3881 4536 3893 4539
rect 3266 4508 3893 4536
rect 3881 4505 3893 4508
rect 3927 4505 3939 4539
rect 5810 4536 5816 4548
rect 3881 4499 3939 4505
rect 3988 4508 5816 4536
rect 3988 4480 4016 4508
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 6029 4539 6087 4545
rect 6029 4505 6041 4539
rect 6075 4536 6087 4539
rect 7834 4536 7840 4548
rect 6075 4508 7840 4536
rect 6075 4505 6087 4508
rect 6029 4499 6087 4505
rect 7834 4496 7840 4508
rect 7892 4496 7898 4548
rect 3970 4428 3976 4480
rect 4028 4428 4034 4480
rect 5626 4428 5632 4480
rect 5684 4428 5690 4480
rect 6181 4471 6239 4477
rect 6181 4437 6193 4471
rect 6227 4468 6239 4471
rect 6730 4468 6736 4480
rect 6227 4440 6736 4468
rect 6227 4437 6239 4440
rect 6181 4431 6239 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 1104 4378 9016 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 9016 4378
rect 1104 4304 9016 4326
rect 5537 4267 5595 4273
rect 5537 4233 5549 4267
rect 5583 4264 5595 4267
rect 5829 4267 5887 4273
rect 5829 4264 5841 4267
rect 5583 4236 5841 4264
rect 5583 4233 5595 4236
rect 5537 4227 5595 4233
rect 5829 4233 5841 4236
rect 5875 4233 5887 4267
rect 5829 4227 5887 4233
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6420 4236 7512 4264
rect 6420 4224 6426 4236
rect 3881 4199 3939 4205
rect 3881 4196 3893 4199
rect 2148 4168 3893 4196
rect 2041 3995 2099 4001
rect 2041 3961 2053 3995
rect 2087 3992 2099 3995
rect 2148 3992 2176 4168
rect 3881 4165 3893 4168
rect 3927 4196 3939 4199
rect 3970 4196 3976 4208
rect 3927 4168 3976 4196
rect 3927 4165 3939 4168
rect 3881 4159 3939 4165
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 4097 4199 4155 4205
rect 4097 4165 4109 4199
rect 4143 4196 4155 4199
rect 4143 4168 4384 4196
rect 4143 4165 4155 4168
rect 4097 4159 4155 4165
rect 4356 4137 4384 4168
rect 4706 4156 4712 4208
rect 4764 4196 4770 4208
rect 5169 4199 5227 4205
rect 4764 4168 5028 4196
rect 4764 4156 4770 4168
rect 5000 4137 5028 4168
rect 5169 4165 5181 4199
rect 5215 4196 5227 4199
rect 5629 4199 5687 4205
rect 5215 4168 5580 4196
rect 5215 4165 5227 4168
rect 5169 4159 5227 4165
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4341 4091 4399 4097
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 4571 4100 4813 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 4801 4091 4859 4097
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5077 4131 5135 4137
rect 5077 4128 5089 4131
rect 5031 4100 5089 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5077 4097 5089 4100
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 2774 4060 2780 4072
rect 2363 4032 2780 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 2774 4020 2780 4032
rect 2832 4060 2838 4072
rect 3510 4060 3516 4072
rect 2832 4032 3516 4060
rect 2832 4020 2838 4032
rect 3510 4020 3516 4032
rect 3568 4020 3574 4072
rect 4816 4060 4844 4091
rect 5184 4060 5212 4159
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5552 4128 5580 4168
rect 5629 4165 5641 4199
rect 5675 4196 5687 4199
rect 5675 4168 5856 4196
rect 5675 4165 5687 4168
rect 5629 4159 5687 4165
rect 5828 4140 5856 4168
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 6822 4196 6828 4208
rect 6512 4168 6828 4196
rect 6512 4156 6518 4168
rect 6822 4156 6828 4168
rect 6880 4196 6886 4208
rect 7484 4205 7512 4236
rect 7009 4199 7067 4205
rect 7009 4196 7021 4199
rect 6880 4168 7021 4196
rect 6880 4156 6886 4168
rect 7009 4165 7021 4168
rect 7055 4165 7067 4199
rect 7009 4159 7067 4165
rect 7469 4199 7527 4205
rect 7469 4165 7481 4199
rect 7515 4165 7527 4199
rect 7469 4159 7527 4165
rect 5552 4100 5672 4128
rect 5353 4091 5411 4097
rect 4816 4032 5212 4060
rect 5368 4060 5396 4091
rect 5534 4060 5540 4072
rect 5368 4032 5540 4060
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5644 4060 5672 4100
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 7742 4128 7748 4140
rect 7699 4100 7748 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 7834 4088 7840 4140
rect 7892 4088 7898 4140
rect 8202 4137 8208 4140
rect 8197 4128 8208 4137
rect 7944 4100 8208 4128
rect 6270 4060 6276 4072
rect 5644 4032 6276 4060
rect 6270 4020 6276 4032
rect 6328 4020 6334 4072
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7944 4060 7972 4100
rect 8197 4091 8208 4100
rect 8202 4088 8208 4091
rect 8260 4088 8266 4140
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 7064 4032 7972 4060
rect 7064 4020 7070 4032
rect 4893 3995 4951 4001
rect 4893 3992 4905 3995
rect 2087 3964 2176 3992
rect 4080 3964 4905 3992
rect 2087 3961 2099 3964
rect 2041 3955 2099 3961
rect 1854 3884 1860 3936
rect 1912 3884 1918 3936
rect 4080 3933 4108 3964
rect 4893 3961 4905 3964
rect 4939 3961 4951 3995
rect 4893 3955 4951 3961
rect 4065 3927 4123 3933
rect 4065 3893 4077 3927
rect 4111 3893 4123 3927
rect 4065 3887 4123 3893
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 4706 3924 4712 3936
rect 4295 3896 4712 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5813 3927 5871 3933
rect 5813 3924 5825 3927
rect 5684 3896 5825 3924
rect 5684 3884 5690 3896
rect 5813 3893 5825 3896
rect 5859 3893 5871 3927
rect 5813 3887 5871 3893
rect 5902 3884 5908 3936
rect 5960 3924 5966 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5960 3896 6009 3924
rect 5960 3884 5966 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 5997 3887 6055 3893
rect 1104 3834 9016 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 9016 3834
rect 1104 3760 9016 3782
rect 1854 3680 1860 3732
rect 1912 3720 1918 3732
rect 2022 3723 2080 3729
rect 2022 3720 2034 3723
rect 1912 3692 2034 3720
rect 1912 3680 1918 3692
rect 2022 3689 2034 3692
rect 2068 3689 2080 3723
rect 2022 3683 2080 3689
rect 3510 3680 3516 3732
rect 3568 3680 3574 3732
rect 5905 3723 5963 3729
rect 5905 3689 5917 3723
rect 5951 3720 5963 3723
rect 6270 3720 6276 3732
rect 5951 3692 6276 3720
rect 5951 3689 5963 3692
rect 5905 3683 5963 3689
rect 6270 3680 6276 3692
rect 6328 3680 6334 3732
rect 7742 3680 7748 3732
rect 7800 3720 7806 3732
rect 8205 3723 8263 3729
rect 8205 3720 8217 3723
rect 7800 3692 8217 3720
rect 7800 3680 7806 3692
rect 8205 3689 8217 3692
rect 8251 3689 8263 3723
rect 8205 3683 8263 3689
rect 1762 3544 1768 3596
rect 1820 3584 1826 3596
rect 4157 3587 4215 3593
rect 4157 3584 4169 3587
rect 1820 3556 4169 3584
rect 1820 3544 1826 3556
rect 4157 3553 4169 3556
rect 4203 3584 4215 3587
rect 4522 3584 4528 3596
rect 4203 3556 4528 3584
rect 4203 3553 4215 3556
rect 4157 3547 4215 3553
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 6730 3544 6736 3596
rect 6788 3544 6794 3596
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3752 3488 3985 3516
rect 3752 3476 3758 3488
rect 3973 3485 3985 3488
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3485 6331 3519
rect 6273 3479 6331 3485
rect 3881 3451 3939 3457
rect 3881 3448 3893 3451
rect 3266 3420 3893 3448
rect 3881 3417 3893 3420
rect 3927 3417 3939 3451
rect 3881 3411 3939 3417
rect 3988 3380 4016 3479
rect 4433 3451 4491 3457
rect 4433 3417 4445 3451
rect 4479 3448 4491 3451
rect 4706 3448 4712 3460
rect 4479 3420 4712 3448
rect 4479 3417 4491 3420
rect 4433 3411 4491 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 6181 3451 6239 3457
rect 6181 3448 6193 3451
rect 5658 3420 6193 3448
rect 6181 3417 6193 3420
rect 6227 3417 6239 3451
rect 6181 3411 6239 3417
rect 6288 3448 6316 3479
rect 6454 3476 6460 3528
rect 6512 3476 6518 3528
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8297 3519 8355 3525
rect 8297 3516 8309 3519
rect 8260 3488 8309 3516
rect 8260 3476 8266 3488
rect 8297 3485 8309 3488
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 7006 3448 7012 3460
rect 6288 3420 7012 3448
rect 6288 3380 6316 3420
rect 7006 3408 7012 3420
rect 7064 3408 7070 3460
rect 8389 3451 8447 3457
rect 8389 3448 8401 3451
rect 7958 3420 8401 3448
rect 8389 3417 8401 3420
rect 8435 3417 8447 3451
rect 8389 3411 8447 3417
rect 3988 3352 6316 3380
rect 1104 3290 9016 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 9016 3290
rect 1104 3216 9016 3238
rect 4433 3179 4491 3185
rect 4433 3145 4445 3179
rect 4479 3176 4491 3179
rect 5534 3176 5540 3188
rect 4479 3148 5540 3176
rect 4479 3145 4491 3148
rect 4433 3139 4491 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 6457 3179 6515 3185
rect 6457 3176 6469 3179
rect 5644 3148 6469 3176
rect 5644 3108 5672 3148
rect 6457 3145 6469 3148
rect 6503 3145 6515 3179
rect 6457 3139 6515 3145
rect 5474 3080 5672 3108
rect 5902 3068 5908 3120
rect 5960 3068 5966 3120
rect 6181 3043 6239 3049
rect 6181 3009 6193 3043
rect 6227 3040 6239 3043
rect 6454 3040 6460 3052
rect 6227 3012 6460 3040
rect 6227 3009 6239 3012
rect 6181 3003 6239 3009
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6549 3043 6607 3049
rect 6549 3009 6561 3043
rect 6595 3040 6607 3043
rect 7006 3040 7012 3052
rect 6595 3012 7012 3040
rect 6595 3009 6607 3012
rect 6549 3003 6607 3009
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 8662 3000 8668 3052
rect 8720 3000 8726 3052
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2836 8079 2839
rect 8570 2836 8576 2848
rect 8067 2808 8576 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 1104 2746 9016 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 9016 2746
rect 1104 2672 9016 2694
rect 8294 2592 8300 2644
rect 8352 2592 8358 2644
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 1104 2202 9016 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 9016 2202
rect 1104 2128 9016 2150
<< via1 >>
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5264 9664 5316 9716
rect 3240 9596 3292 9648
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 3424 9392 3476 9444
rect 3976 9392 4028 9444
rect 5816 9528 5868 9580
rect 6460 9528 6512 9580
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 5632 9392 5684 9444
rect 3608 9324 3660 9376
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 5724 9324 5776 9376
rect 6644 9324 6696 9376
rect 7012 9324 7064 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2228 9163 2280 9172
rect 2228 9129 2237 9163
rect 2237 9129 2271 9163
rect 2271 9129 2280 9163
rect 2228 9120 2280 9129
rect 5632 9120 5684 9172
rect 3148 9095 3200 9104
rect 3148 9061 3157 9095
rect 3157 9061 3191 9095
rect 3191 9061 3200 9095
rect 3148 9052 3200 9061
rect 2596 8984 2648 9036
rect 848 8916 900 8968
rect 3608 8984 3660 9036
rect 7012 9095 7064 9104
rect 7012 9061 7021 9095
rect 7021 9061 7055 9095
rect 7055 9061 7064 9095
rect 7012 9052 7064 9061
rect 2872 8891 2924 8900
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 2872 8857 2881 8891
rect 2881 8857 2915 8891
rect 2915 8857 2924 8891
rect 2872 8848 2924 8857
rect 3240 8780 3292 8832
rect 5724 8984 5776 9036
rect 3976 8959 4028 8968
rect 3976 8925 3985 8959
rect 3985 8925 4019 8959
rect 4019 8925 4028 8959
rect 3976 8916 4028 8925
rect 4804 8959 4856 8968
rect 4804 8925 4813 8959
rect 4813 8925 4847 8959
rect 4847 8925 4856 8959
rect 4804 8916 4856 8925
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 6828 8984 6880 9036
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 4252 8780 4304 8832
rect 5448 8780 5500 8832
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 8116 8916 8168 8968
rect 7196 8823 7248 8832
rect 7196 8789 7205 8823
rect 7205 8789 7239 8823
rect 7239 8789 7248 8823
rect 7196 8780 7248 8789
rect 8208 8780 8260 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2412 8619 2464 8628
rect 2412 8585 2421 8619
rect 2421 8585 2455 8619
rect 2455 8585 2464 8619
rect 2412 8576 2464 8585
rect 2504 8576 2556 8628
rect 3332 8576 3384 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2136 8347 2188 8356
rect 2136 8313 2145 8347
rect 2145 8313 2179 8347
rect 2179 8313 2188 8347
rect 2136 8304 2188 8313
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 2596 8483 2648 8492
rect 2596 8449 2605 8483
rect 2605 8449 2639 8483
rect 2639 8449 2648 8483
rect 2596 8440 2648 8449
rect 2964 8440 3016 8492
rect 3240 8440 3292 8492
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 4252 8576 4304 8628
rect 3792 8483 3844 8492
rect 3792 8449 3801 8483
rect 3801 8449 3835 8483
rect 3835 8449 3844 8483
rect 3792 8440 3844 8449
rect 5448 8551 5500 8560
rect 5448 8517 5457 8551
rect 5457 8517 5491 8551
rect 5491 8517 5500 8551
rect 5448 8508 5500 8517
rect 4252 8483 4304 8492
rect 4252 8449 4261 8483
rect 4261 8449 4295 8483
rect 4295 8449 4304 8483
rect 4252 8440 4304 8449
rect 4344 8440 4396 8492
rect 4528 8440 4580 8492
rect 5632 8440 5684 8492
rect 6184 8508 6236 8560
rect 6276 8440 6328 8492
rect 1492 8236 1544 8288
rect 2596 8236 2648 8288
rect 2780 8279 2832 8288
rect 2780 8245 2789 8279
rect 2789 8245 2823 8279
rect 2823 8245 2832 8279
rect 2780 8236 2832 8245
rect 3516 8236 3568 8288
rect 4068 8304 4120 8356
rect 4804 8304 4856 8356
rect 5448 8304 5500 8356
rect 6460 8440 6512 8492
rect 7748 8415 7800 8424
rect 7748 8381 7757 8415
rect 7757 8381 7791 8415
rect 7791 8381 7800 8415
rect 7748 8372 7800 8381
rect 8024 8415 8076 8424
rect 8024 8381 8033 8415
rect 8033 8381 8067 8415
rect 8067 8381 8076 8415
rect 8024 8372 8076 8381
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8392 8372 8444 8424
rect 6552 8304 6604 8356
rect 6920 8279 6972 8288
rect 6920 8245 6929 8279
rect 6929 8245 6963 8279
rect 6963 8245 6972 8279
rect 6920 8236 6972 8245
rect 7472 8347 7524 8356
rect 7472 8313 7481 8347
rect 7481 8313 7515 8347
rect 7515 8313 7524 8347
rect 7472 8304 7524 8313
rect 7564 8236 7616 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 1860 8032 1912 8084
rect 7748 8075 7800 8084
rect 7748 8041 7757 8075
rect 7757 8041 7791 8075
rect 7791 8041 7800 8075
rect 7748 8032 7800 8041
rect 8392 8075 8444 8084
rect 8392 8041 8401 8075
rect 8401 8041 8435 8075
rect 8435 8041 8444 8075
rect 8392 8032 8444 8041
rect 848 7828 900 7880
rect 1860 7828 1912 7880
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 6920 7896 6972 7948
rect 2964 7828 3016 7880
rect 3148 7828 3200 7880
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 6184 7828 6236 7880
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 7288 7871 7340 7880
rect 7288 7837 7297 7871
rect 7297 7837 7331 7871
rect 7331 7837 7340 7871
rect 7288 7828 7340 7837
rect 7564 7871 7616 7880
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 8024 7896 8076 7948
rect 6552 7760 6604 7812
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8576 7760 8628 7812
rect 2872 7692 2924 7744
rect 5908 7692 5960 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1860 7531 1912 7540
rect 1860 7497 1869 7531
rect 1869 7497 1903 7531
rect 1903 7497 1912 7531
rect 1860 7488 1912 7497
rect 2596 7488 2648 7540
rect 3424 7488 3476 7540
rect 1768 7420 1820 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 2688 7352 2740 7404
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3424 7395 3476 7404
rect 3424 7361 3431 7395
rect 3431 7361 3476 7395
rect 3424 7352 3476 7361
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 3608 7284 3660 7336
rect 4528 7352 4580 7404
rect 5816 7420 5868 7472
rect 4436 7327 4488 7336
rect 4436 7293 4445 7327
rect 4445 7293 4479 7327
rect 4479 7293 4488 7327
rect 4436 7284 4488 7293
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6644 7352 6696 7404
rect 8116 7352 8168 7404
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 5448 7216 5500 7268
rect 5540 7216 5592 7268
rect 6276 7284 6328 7336
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 2780 7148 2832 7200
rect 3516 7148 3568 7200
rect 4068 7148 4120 7200
rect 4436 7148 4488 7200
rect 6368 7148 6420 7200
rect 6736 7148 6788 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3148 6987 3200 6996
rect 3148 6953 3157 6987
rect 3157 6953 3191 6987
rect 3191 6953 3200 6987
rect 3148 6944 3200 6953
rect 2688 6876 2740 6928
rect 3608 6876 3660 6928
rect 6184 6876 6236 6928
rect 6552 6876 6604 6928
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 1768 6783 1820 6792
rect 1768 6749 1777 6783
rect 1777 6749 1811 6783
rect 1811 6749 1820 6783
rect 1768 6740 1820 6749
rect 2964 6740 3016 6792
rect 5264 6740 5316 6792
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 5908 6740 5960 6792
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 2780 6672 2832 6724
rect 6184 6715 6236 6724
rect 6184 6681 6193 6715
rect 6193 6681 6227 6715
rect 6227 6681 6236 6715
rect 6184 6672 6236 6681
rect 1952 6647 2004 6656
rect 1952 6613 1961 6647
rect 1961 6613 1995 6647
rect 1995 6613 2004 6647
rect 1952 6604 2004 6613
rect 5632 6604 5684 6656
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 7196 6808 7248 6860
rect 7104 6715 7156 6724
rect 7104 6681 7113 6715
rect 7113 6681 7147 6715
rect 7147 6681 7156 6715
rect 7104 6672 7156 6681
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 8208 6783 8260 6792
rect 8208 6749 8217 6783
rect 8217 6749 8251 6783
rect 8251 6749 8260 6783
rect 8208 6740 8260 6749
rect 7840 6715 7892 6724
rect 7840 6681 7849 6715
rect 7849 6681 7883 6715
rect 7883 6681 7892 6715
rect 7840 6672 7892 6681
rect 8300 6647 8352 6656
rect 8300 6613 8309 6647
rect 8309 6613 8343 6647
rect 8343 6613 8352 6647
rect 8300 6604 8352 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2780 6400 2832 6452
rect 1768 6375 1820 6384
rect 1768 6341 1777 6375
rect 1777 6341 1811 6375
rect 1811 6341 1820 6375
rect 1768 6332 1820 6341
rect 3148 6332 3200 6384
rect 3608 6443 3660 6452
rect 3608 6409 3617 6443
rect 3617 6409 3651 6443
rect 3651 6409 3660 6443
rect 3608 6400 3660 6409
rect 4068 6443 4120 6452
rect 4068 6409 4077 6443
rect 4077 6409 4111 6443
rect 4111 6409 4120 6443
rect 4068 6400 4120 6409
rect 4620 6400 4672 6452
rect 4896 6400 4948 6452
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 4068 6264 4120 6316
rect 7196 6375 7248 6384
rect 7196 6341 7205 6375
rect 7205 6341 7239 6375
rect 7239 6341 7248 6375
rect 7196 6332 7248 6341
rect 8300 6264 8352 6316
rect 1768 6128 1820 6180
rect 4068 6128 4120 6180
rect 4896 6239 4948 6248
rect 4896 6205 4905 6239
rect 4905 6205 4939 6239
rect 4939 6205 4948 6239
rect 4896 6196 4948 6205
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 6920 6196 6972 6205
rect 2228 6060 2280 6112
rect 4712 6060 4764 6112
rect 7932 6060 7984 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 1492 5856 1544 5908
rect 2136 5788 2188 5840
rect 1952 5720 2004 5772
rect 1584 5516 1636 5568
rect 2228 5627 2280 5636
rect 2228 5593 2253 5627
rect 2253 5593 2280 5627
rect 3148 5899 3200 5908
rect 3148 5865 3157 5899
rect 3157 5865 3191 5899
rect 3191 5865 3200 5899
rect 3148 5856 3200 5865
rect 4252 5856 4304 5908
rect 4896 5856 4948 5908
rect 5264 5856 5316 5908
rect 7840 5856 7892 5908
rect 8300 5788 8352 5840
rect 4620 5720 4672 5772
rect 3700 5652 3752 5704
rect 7012 5720 7064 5772
rect 8208 5720 8260 5772
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 2228 5584 2280 5593
rect 3884 5584 3936 5636
rect 4068 5584 4120 5636
rect 3516 5516 3568 5568
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 7472 5695 7524 5704
rect 7472 5661 7481 5695
rect 7481 5661 7515 5695
rect 7515 5661 7524 5695
rect 7472 5652 7524 5661
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 7104 5584 7156 5636
rect 7748 5584 7800 5636
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 7196 5559 7248 5568
rect 7196 5525 7205 5559
rect 7205 5525 7239 5559
rect 7239 5525 7248 5559
rect 7196 5516 7248 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 6920 5312 6972 5364
rect 4252 5287 4304 5296
rect 4252 5253 4261 5287
rect 4261 5253 4295 5287
rect 4295 5253 4304 5287
rect 4252 5244 4304 5253
rect 4436 5287 4488 5296
rect 4436 5253 4445 5287
rect 4445 5253 4479 5287
rect 4479 5253 4488 5287
rect 4436 5244 4488 5253
rect 1492 5219 1544 5228
rect 1492 5185 1501 5219
rect 1501 5185 1535 5219
rect 1535 5185 1544 5219
rect 1492 5176 1544 5185
rect 1584 5219 1636 5228
rect 1584 5185 1593 5219
rect 1593 5185 1627 5219
rect 1627 5185 1636 5219
rect 1584 5176 1636 5185
rect 4712 5176 4764 5228
rect 5540 5176 5592 5228
rect 6184 5176 6236 5228
rect 7196 5244 7248 5296
rect 1768 5108 1820 5160
rect 5816 5108 5868 5160
rect 6276 5040 6328 5092
rect 6828 5151 6880 5160
rect 6828 5117 6837 5151
rect 6837 5117 6871 5151
rect 6871 5117 6880 5151
rect 6828 5108 6880 5117
rect 7472 5108 7524 5160
rect 8300 5108 8352 5160
rect 2044 4972 2096 5024
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 8576 5015 8628 5024
rect 8576 4981 8585 5015
rect 8585 4981 8619 5015
rect 8619 4981 8628 5015
rect 8576 4972 8628 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 3516 4811 3568 4820
rect 3516 4777 3525 4811
rect 3525 4777 3559 4811
rect 3559 4777 3568 4811
rect 3516 4768 3568 4777
rect 6552 4768 6604 4820
rect 7380 4768 7432 4820
rect 6828 4700 6880 4752
rect 2044 4675 2096 4684
rect 2044 4641 2053 4675
rect 2053 4641 2087 4675
rect 2087 4641 2096 4675
rect 2044 4632 2096 4641
rect 6552 4675 6604 4684
rect 6552 4641 6561 4675
rect 6561 4641 6595 4675
rect 6595 4641 6604 4675
rect 6552 4632 6604 4641
rect 1768 4607 1820 4616
rect 1768 4573 1777 4607
rect 1777 4573 1811 4607
rect 1811 4573 1820 4607
rect 1768 4564 1820 4573
rect 3700 4564 3752 4616
rect 6368 4564 6420 4616
rect 8576 4632 8628 4684
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 5816 4539 5868 4548
rect 5816 4505 5825 4539
rect 5825 4505 5859 4539
rect 5859 4505 5868 4539
rect 5816 4496 5868 4505
rect 7840 4496 7892 4548
rect 3976 4428 4028 4480
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 6736 4428 6788 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 6368 4224 6420 4276
rect 3976 4156 4028 4208
rect 4712 4199 4764 4208
rect 4712 4165 4721 4199
rect 4721 4165 4755 4199
rect 4755 4165 4764 4199
rect 4712 4156 4764 4165
rect 2780 4020 2832 4072
rect 3516 4020 3568 4072
rect 6460 4156 6512 4208
rect 6828 4156 6880 4208
rect 5540 4020 5592 4072
rect 5816 4088 5868 4140
rect 7748 4088 7800 4140
rect 7840 4131 7892 4140
rect 7840 4097 7849 4131
rect 7849 4097 7883 4131
rect 7883 4097 7892 4131
rect 7840 4088 7892 4097
rect 8208 4131 8260 4140
rect 6276 4020 6328 4072
rect 7012 4020 7064 4072
rect 8208 4097 8209 4131
rect 8209 4097 8243 4131
rect 8243 4097 8260 4131
rect 8208 4088 8260 4097
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 4712 3884 4764 3936
rect 5632 3884 5684 3936
rect 5908 3884 5960 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 1860 3680 1912 3732
rect 3516 3723 3568 3732
rect 3516 3689 3525 3723
rect 3525 3689 3559 3723
rect 3559 3689 3568 3723
rect 3516 3680 3568 3689
rect 6276 3680 6328 3732
rect 7748 3680 7800 3732
rect 1768 3587 1820 3596
rect 1768 3553 1777 3587
rect 1777 3553 1811 3587
rect 1811 3553 1820 3587
rect 1768 3544 1820 3553
rect 4528 3544 4580 3596
rect 6736 3587 6788 3596
rect 6736 3553 6745 3587
rect 6745 3553 6779 3587
rect 6779 3553 6788 3587
rect 6736 3544 6788 3553
rect 3700 3476 3752 3528
rect 4712 3408 4764 3460
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 8208 3476 8260 3528
rect 7012 3408 7064 3460
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5540 3136 5592 3188
rect 5908 3111 5960 3120
rect 5908 3077 5917 3111
rect 5917 3077 5951 3111
rect 5951 3077 5960 3111
rect 5908 3068 5960 3077
rect 6460 3000 6512 3052
rect 7012 3000 7064 3052
rect 8668 3043 8720 3052
rect 8668 3009 8677 3043
rect 8677 3009 8711 3043
rect 8711 3009 8720 3043
rect 8668 3000 8720 3009
rect 8576 2796 8628 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 8300 2635 8352 2644
rect 8300 2601 8309 2635
rect 8309 2601 8343 2635
rect 8343 2601 8352 2635
rect 8300 2592 8352 2601
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 3238 11549 3294 12349
rect 5170 11549 5226 12349
rect 5814 11549 5870 12349
rect 6458 11549 6514 12349
rect 3252 9654 3280 11549
rect 5184 10010 5212 11549
rect 5184 9982 5304 10010
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9722 5304 9982
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 5828 9586 5856 11549
rect 6472 9586 6500 11549
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 846 9072 902 9081
rect 2240 9058 2268 9114
rect 3148 9104 3200 9110
rect 2240 9042 2636 9058
rect 3148 9046 3200 9052
rect 2240 9036 2648 9042
rect 2240 9030 2596 9036
rect 846 9007 902 9016
rect 860 8974 888 9007
rect 2596 8978 2648 8984
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2424 8634 2452 8774
rect 2516 8634 2544 8774
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2516 8498 2544 8570
rect 2608 8498 2636 8978
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2596 8492 2648 8498
rect 2884 8480 2912 8842
rect 2964 8492 3016 8498
rect 2884 8452 2964 8480
rect 2596 8434 2648 8440
rect 2964 8434 3016 8440
rect 1412 8265 1440 8434
rect 1492 8288 1544 8294
rect 1398 8256 1454 8265
rect 1492 8230 1544 8236
rect 1398 8191 1454 8200
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 1504 7410 1532 8230
rect 1872 8090 1900 8434
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1872 7546 1900 7822
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1768 7472 1820 7478
rect 1768 7414 1820 7420
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1780 6798 1808 7414
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1780 6390 1808 6734
rect 1964 6662 1992 8434
rect 2134 8392 2190 8401
rect 2134 8327 2136 8336
rect 2188 8327 2190 8336
rect 2136 8298 2188 8304
rect 2608 8294 2636 8434
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2780 8288 2832 8294
rect 2780 8230 2832 8236
rect 2792 7954 2820 8230
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2976 7886 3004 8434
rect 3160 7886 3188 9046
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8498 3280 8774
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3344 8498 3372 8570
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2608 7546 2636 7822
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2884 7410 2912 7686
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 2700 6934 2728 7346
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2688 6928 2740 6934
rect 2688 6870 2740 6876
rect 2792 6730 2820 7142
rect 2976 6798 3004 7822
rect 3436 7546 3464 9386
rect 3620 9382 3648 9522
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 3976 9444 4028 9450
rect 3976 9386 4028 9392
rect 3608 9376 3660 9382
rect 3608 9318 3660 9324
rect 3620 9042 3648 9318
rect 3608 9036 3660 9042
rect 3608 8978 3660 8984
rect 3988 8974 4016 9386
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 5368 8974 5396 9318
rect 5552 8974 5580 9454
rect 5632 9444 5684 9450
rect 5632 9386 5684 9392
rect 5644 9178 5672 9386
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4264 8634 4292 8774
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4264 8498 4292 8570
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3792 8492 3844 8498
rect 4252 8492 4304 8498
rect 3844 8452 4200 8480
rect 3792 8434 3844 8440
rect 3528 8294 3556 8434
rect 4066 8392 4122 8401
rect 4172 8378 4200 8452
rect 4252 8434 4304 8440
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4528 8492 4580 8498
rect 4580 8452 4660 8480
rect 4528 8434 4580 8440
rect 4356 8378 4384 8434
rect 4172 8350 4384 8378
rect 4066 8327 4068 8336
rect 4120 8327 4122 8336
rect 4068 8298 4120 8304
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3436 7410 3464 7482
rect 3528 7410 3556 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 4528 7404 4580 7410
rect 4632 7392 4660 8452
rect 4816 8362 4844 8910
rect 5448 8832 5500 8838
rect 5448 8774 5500 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5460 8566 5488 8774
rect 5448 8560 5500 8566
rect 5448 8502 5500 8508
rect 4804 8356 4856 8362
rect 4804 8298 4856 8304
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4580 7364 4660 7392
rect 4528 7346 4580 7352
rect 3160 7002 3188 7346
rect 3528 7206 3556 7346
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 3516 7200 3568 7206
rect 3516 7142 3568 7148
rect 3148 6996 3200 7002
rect 3148 6938 3200 6944
rect 2964 6792 3016 6798
rect 2964 6734 3016 6740
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1768 6384 1820 6390
rect 1768 6326 1820 6332
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1504 5234 1532 5850
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1596 5234 1624 5510
rect 1492 5228 1544 5234
rect 1492 5170 1544 5176
rect 1584 5228 1636 5234
rect 1584 5170 1636 5176
rect 1780 5166 1808 6122
rect 1964 5778 1992 6598
rect 2792 6458 2820 6666
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2148 5846 2176 6190
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2136 5840 2188 5846
rect 2136 5782 2188 5788
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 2240 5642 2268 6054
rect 2228 5636 2280 5642
rect 2228 5578 2280 5584
rect 1768 5160 1820 5166
rect 1768 5102 1820 5108
rect 1780 4622 1808 5102
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2056 4690 2084 4966
rect 2044 4684 2096 4690
rect 2044 4626 2096 4632
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1780 3602 1808 4558
rect 2792 4078 2820 6394
rect 3148 6384 3200 6390
rect 3148 6326 3200 6332
rect 3160 5914 3188 6326
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3528 5574 3556 7142
rect 3620 6934 3648 7278
rect 4448 7206 4476 7278
rect 4068 7200 4120 7206
rect 4068 7142 4120 7148
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 3608 6928 3660 6934
rect 3608 6870 3660 6876
rect 3620 6458 3648 6870
rect 4080 6458 4108 7142
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4632 6458 4660 7364
rect 5460 7274 5488 8298
rect 5552 7886 5580 8910
rect 5644 8498 5672 9114
rect 5736 9042 5764 9318
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 6656 8974 6684 9318
rect 6840 9042 6868 9522
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 7024 9110 7052 9318
rect 7012 9104 7064 9110
rect 7012 9046 7064 9052
rect 6828 9036 6880 9042
rect 6828 8978 6880 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6196 8566 6224 8774
rect 6184 8560 6236 8566
rect 6184 8502 6236 8508
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 6196 7886 6224 8502
rect 6276 8492 6328 8498
rect 6460 8492 6512 8498
rect 6328 8452 6460 8480
rect 6276 8434 6328 8440
rect 6460 8434 6512 8440
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5540 7268 5592 7274
rect 5540 7210 5592 7216
rect 5460 6798 5488 7210
rect 5552 6798 5580 7210
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4080 6322 4108 6394
rect 4068 6316 4120 6322
rect 4068 6258 4120 6264
rect 4908 6254 4936 6394
rect 4896 6248 4948 6254
rect 4896 6190 4948 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3516 5568 3568 5574
rect 3516 5510 3568 5516
rect 3528 4826 3556 5510
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3712 4622 3740 5646
rect 4080 5642 4108 6122
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3896 5522 3924 5578
rect 3896 5494 4016 5522
rect 3700 4616 3752 4622
rect 3700 4558 3752 4564
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 3516 4072 3568 4078
rect 3516 4014 3568 4020
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1872 3738 1900 3878
rect 3528 3738 3556 4014
rect 1860 3732 1912 3738
rect 1860 3674 1912 3680
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 1768 3596 1820 3602
rect 1768 3538 1820 3544
rect 3712 3534 3740 4558
rect 3988 4486 4016 5494
rect 4264 5302 4292 5850
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4434 5536 4490 5545
rect 4434 5471 4490 5480
rect 4448 5302 4476 5471
rect 4252 5296 4304 5302
rect 4252 5238 4304 5244
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3988 4214 4016 4422
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3618 4660 5714
rect 4724 5234 4752 6054
rect 4908 5914 4936 6190
rect 5276 5914 5304 6734
rect 5644 6662 5672 7278
rect 5828 6866 5856 7414
rect 5920 7410 5948 7686
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5920 6798 5948 7346
rect 6288 7342 6316 8434
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 7818 6592 8298
rect 6552 7812 6604 7818
rect 6552 7754 6604 7760
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6184 6928 6236 6934
rect 6184 6870 6236 6876
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 6196 6730 6224 6870
rect 6184 6724 6236 6730
rect 6184 6666 6236 6672
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 6196 5234 6224 6666
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 4724 4214 4752 5170
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 5552 4078 5580 5170
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4554 5856 5102
rect 6288 5098 6316 7278
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6380 6798 6408 7142
rect 6564 6934 6592 7754
rect 6656 7410 6684 8910
rect 7196 8832 7248 8838
rect 7196 8774 7248 8780
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 7954 6960 8230
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 7208 7886 7236 8774
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7288 7880 7340 7886
rect 7288 7822 7340 7828
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6552 6928 6604 6934
rect 6552 6870 6604 6876
rect 6748 6798 6776 7142
rect 7300 7018 7328 7822
rect 7116 6990 7328 7018
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 7116 6730 7144 6990
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7104 6724 7156 6730
rect 7104 6666 7156 6672
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6276 5092 6328 5098
rect 6276 5034 6328 5040
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4540 3602 4660 3618
rect 4528 3596 4660 3602
rect 4580 3590 4660 3596
rect 4528 3538 4580 3544
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 4724 3466 4752 3878
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5552 3194 5580 4014
rect 5644 3942 5672 4422
rect 5828 4146 5856 4490
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 6288 4078 6316 5034
rect 6380 5030 6408 5646
rect 6552 5568 6604 5574
rect 6932 5522 6960 6190
rect 7012 5772 7064 5778
rect 7012 5714 7064 5720
rect 6552 5510 6604 5516
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4622 6408 4966
rect 6564 4826 6592 5510
rect 6840 5494 6960 5522
rect 6840 5166 6868 5494
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6828 5160 6880 5166
rect 6828 5102 6880 5108
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6564 4690 6592 4762
rect 6840 4758 6868 5102
rect 6828 4752 6880 4758
rect 6828 4694 6880 4700
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6380 4282 6408 4558
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5920 3126 5948 3878
rect 6288 3738 6316 4014
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6472 3534 6500 4150
rect 6748 3602 6776 4422
rect 6840 4214 6868 4694
rect 6932 4622 6960 5306
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 7024 4078 7052 5714
rect 7116 5642 7144 6666
rect 7208 6390 7236 6802
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7484 5710 7512 8298
rect 7564 8288 7616 8294
rect 7564 8230 7616 8236
rect 7576 7886 7604 8230
rect 7760 8090 7788 8366
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 8036 7954 8064 8366
rect 8024 7948 8076 7954
rect 8024 7890 8076 7896
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 8128 7410 8156 8910
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8498 8248 8774
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 7886 8248 8434
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8404 8090 8432 8366
rect 8392 8084 8444 8090
rect 8392 8026 8444 8032
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8128 6798 8156 7346
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7852 5914 7880 6666
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7944 5710 7972 6054
rect 8220 5778 8248 6734
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8312 6322 8340 6598
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 7104 5636 7156 5642
rect 7104 5578 7156 5584
rect 7196 5568 7248 5574
rect 7196 5510 7248 5516
rect 7208 5302 7236 5510
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7392 4826 7420 5646
rect 7484 5166 7512 5646
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7380 4820 7432 4826
rect 7380 4762 7432 4768
rect 7760 4146 7788 5578
rect 8312 5545 8340 5782
rect 8588 5710 8616 7754
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8680 6905 8708 7278
rect 8666 6896 8722 6905
rect 8666 6831 8722 6840
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8298 5536 8354 5545
rect 8298 5471 8354 5480
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7852 4146 7880 4490
rect 8312 4146 8340 5102
rect 8588 5030 8616 5646
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4690 8616 4966
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 6472 3058 6500 3470
rect 7024 3466 7052 4014
rect 7760 3738 7788 4082
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 8220 3534 8248 4082
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8666 3496 8722 3505
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 7024 3058 7052 3402
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 8220 2774 8248 3470
rect 8666 3431 8722 3440
rect 8680 3058 8708 3431
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 8220 2746 8340 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 8312 2650 8340 2746
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8588 2446 8616 2790
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
<< via2 >>
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 846 9016 902 9072
rect 1398 8200 1454 8256
rect 846 7656 902 7712
rect 2134 8356 2190 8392
rect 2134 8336 2136 8356
rect 2136 8336 2188 8356
rect 2188 8336 2190 8356
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4066 8356 4122 8392
rect 4066 8336 4068 8356
rect 4068 8336 4120 8356
rect 4120 8336 4122 8356
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4434 5480 4490 5536
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 8666 6840 8722 6896
rect 8298 5480 8354 5536
rect 8666 3440 8722 3496
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 0 8848 800 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 2129 8394 2195 8397
rect 4061 8394 4127 8397
rect 2129 8392 4127 8394
rect 2129 8336 2134 8392
rect 2190 8336 4066 8392
rect 4122 8336 4127 8392
rect 2129 8334 4127 8336
rect 2129 8331 2195 8334
rect 4061 8331 4127 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 0 7488 800 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 8661 6898 8727 6901
rect 9405 6898 10205 6928
rect 8661 6896 10205 6898
rect 8661 6840 8666 6896
rect 8722 6840 10205 6896
rect 8661 6838 10205 6840
rect 8661 6835 8727 6838
rect 9405 6808 10205 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5538 800 5568
rect 4429 5538 4495 5541
rect 0 5536 4495 5538
rect 0 5480 4434 5536
rect 4490 5480 4495 5536
rect 0 5478 4495 5480
rect 0 5448 800 5478
rect 4429 5475 4495 5478
rect 8293 5538 8359 5541
rect 9405 5538 10205 5568
rect 8293 5536 10205 5538
rect 8293 5480 8298 5536
rect 8354 5480 10205 5536
rect 8293 5478 10205 5480
rect 8293 5475 8359 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 9405 5448 10205 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 8661 3498 8727 3501
rect 9405 3498 10205 3528
rect 8661 3496 10205 3498
rect 8661 3440 8666 3496
rect 8722 3440 10205 3496
rect 8661 3438 10205 3440
rect 8661 3435 8727 3438
rect 9405 3408 10205 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 9280 4528 9840
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 9824 5188 9840
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _073_
timestamp 0
transform -1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 0
transform -1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 0
transform 1 0 5520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _076_
timestamp 0
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 0
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _078_
timestamp 0
transform 1 0 3036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _079_
timestamp 0
transform 1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _080_
timestamp 0
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _081_
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _082_
timestamp 0
transform -1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _083_
timestamp 0
transform 1 0 2024 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _084_
timestamp 0
transform 1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _085_
timestamp 0
transform 1 0 5336 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _086_
timestamp 0
transform -1 0 6716 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _087_
timestamp 0
transform 1 0 7268 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _088_
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _089_
timestamp 0
transform -1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _090_
timestamp 0
transform 1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _091_
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _092_
timestamp 0
transform 1 0 1472 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _093_
timestamp 0
transform 1 0 2300 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _094_
timestamp 0
transform -1 0 2208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _095_
timestamp 0
transform 1 0 3128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _096_
timestamp 0
transform 1 0 4600 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _097_
timestamp 0
transform -1 0 5520 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _098_
timestamp 0
transform 1 0 3864 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _099_
timestamp 0
transform 1 0 5244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _100_
timestamp 0
transform 1 0 5796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _101_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _102_
timestamp 0
transform 1 0 6440 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _103_
timestamp 0
transform 1 0 6808 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _104_
timestamp 0
transform 1 0 6716 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _105_
timestamp 0
transform 1 0 6992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _106_
timestamp 0
transform 1 0 7820 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_4  _107_
timestamp 0
transform -1 0 8740 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _108_
timestamp 0
transform -1 0 2392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _109_
timestamp 0
transform -1 0 1840 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _110_
timestamp 0
transform 1 0 2024 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _111_
timestamp 0
transform -1 0 2024 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _112_
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _113_
timestamp 0
transform 1 0 3772 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 0
transform -1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _115_
timestamp 0
transform 1 0 4416 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _116_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _117_
timestamp 0
transform -1 0 5060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _118_
timestamp 0
transform -1 0 4784 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _119_
timestamp 0
transform 1 0 3864 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _120_
timestamp 0
transform -1 0 6808 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 0
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _122_
timestamp 0
transform -1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _123_
timestamp 0
transform 1 0 5612 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _124_
timestamp 0
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _125_
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _126_
timestamp 0
transform 1 0 5796 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _127_
timestamp 0
transform 1 0 6256 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _128_
timestamp 0
transform -1 0 7636 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _129_
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _130_
timestamp 0
transform -1 0 6256 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _131_
timestamp 0
transform 1 0 2576 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _132_
timestamp 0
transform 1 0 3220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _133_
timestamp 0
transform 1 0 4048 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _134_
timestamp 0
transform -1 0 5796 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _135_
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _136_
timestamp 0
transform 1 0 6348 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _137_
timestamp 0
transform -1 0 7912 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 0
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 0
transform -1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 0
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 0
transform -1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 0
transform -1 0 6348 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 0
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 0
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 0
transform 1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _146_
timestamp 0
transform 1 0 6900 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _147_
timestamp 0
transform 1 0 1748 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _148_
timestamp 0
transform 1 0 1840 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _149_
timestamp 0
transform 1 0 1748 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _150_
timestamp 0
transform 1 0 4232 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _151_
timestamp 0
transform 1 0 4140 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _152_
timestamp 0
transform -1 0 6256 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _153_
timestamp 0
transform 1 0 6440 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _154_
timestamp 0
transform 1 0 6808 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform -1 0 3680 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform 1 0 6900 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 0
transform 1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp 0
transform 1 0 4324 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_60
timestamp 0
transform 1 0 6624 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp 0
transform 1 0 7728 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_32
timestamp 0
transform 1 0 4048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 0
transform 1 0 6348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_81
timestamp 0
transform 1 0 8556 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_7
timestamp 0
transform 1 0 1748 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_14
timestamp 0
transform 1 0 2392 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_26
timestamp 0
transform 1 0 3496 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 0
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_74
timestamp 0
transform 1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_80
timestamp 0
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_32
timestamp 0
transform 1 0 4048 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 0
transform 1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 0
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_32
timestamp 0
transform 1 0 4048 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 0
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_60
timestamp 0
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_43
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_10
timestamp 0
transform 1 0 2024 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_18
timestamp 0
transform 1 0 2760 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 0
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 0
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_80
timestamp 0
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_12
timestamp 0
transform 1 0 2208 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_31
timestamp 0
transform 1 0 3956 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 0
transform 1 0 4876 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp 0
transform 1 0 5244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_62
timestamp 0
transform 1 0 6808 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_70
timestamp 0
transform 1 0 7544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_20
timestamp 0
transform 1 0 2944 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 0
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_47
timestamp 0
transform 1 0 5428 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_51
timestamp 0
transform 1 0 5796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_57
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_63
timestamp 0
transform 1 0 6900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_80
timestamp 0
transform 1 0 8464 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_19
timestamp 0
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_64
timestamp 0
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_36
timestamp 0
transform 1 0 4416 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_45
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_80
timestamp 0
transform 1 0 8464 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 0
transform 1 0 3220 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_32
timestamp 0
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_44
timestamp 0
transform 1 0 5152 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_65
timestamp 0
transform 1 0 7084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_77
timestamp 0
transform 1 0 8188 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 8740 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 8740 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform 1 0 3772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform -1 0 6164 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 0
transform -1 0 8740 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp 0
transform -1 0 8740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 0
transform -1 0 8004 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_14
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_15
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_16
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 9016 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_17
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_18
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 9016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_19
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 9016 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_20
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_21
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 9016 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_22
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 9016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_23
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 9016 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_24
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 9016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_25
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 9016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_26
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 9016 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_27
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 9016 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_30
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_31
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_32
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_33
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_34
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_35
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_36
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_37
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_38
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_39
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_40
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_41
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_42
timestamp 0
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_43
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
<< labels >>
rlabel metal1 s 5060 9792 5060 9792 4 VGND
rlabel metal1 s 5060 9248 5060 9248 4 VPWR
rlabel metal1 s 1968 3706 1968 3706 4 _000_
rlabel metal1 s 2300 5814 2300 5814 4 _001_
rlabel metal2 s 2070 4828 2070 4828 4 _002_
rlabel metal1 s 4370 5610 4370 5610 4 _003_
rlabel metal1 s 4600 3434 4600 3434 4 _004_
rlabel metal2 s 5934 3502 5934 3502 4 _005_
rlabel metal2 s 6762 4012 6762 4012 4 _006_
rlabel metal1 s 7176 5270 7176 5270 4 _007_
rlabel metal1 s 7507 6834 7507 6834 4 _008_
rlabel metal2 s 8326 6460 8326 6460 4 _009_
rlabel metal1 s 3595 3434 3595 3434 4 _010_
rlabel metal2 s 3174 6120 3174 6120 4 _011_
rlabel metal1 s 3595 4522 3595 4522 4 _012_
rlabel metal1 s 5987 5610 5987 5610 4 _013_
rlabel metal1 s 5941 3434 5941 3434 4 _014_
rlabel metal1 s 6072 3162 6072 3162 4 _015_
rlabel metal1 s 8195 3434 8195 3434 4 _016_
rlabel metal2 s 8326 4624 8326 4624 4 _017_
rlabel metal1 s 7498 6698 7498 6698 4 _018_
rlabel metal2 s 6762 6970 6762 6970 4 _019_
rlabel metal2 s 5934 7548 5934 7548 4 _020_
rlabel metal1 s 4370 7276 4370 7276 4 _021_
rlabel metal2 s 4002 9180 4002 9180 4 _022_
rlabel metal2 s 2898 7548 2898 7548 4 _023_
rlabel metal2 s 3174 7174 3174 7174 4 _024_
rlabel metal1 s 2346 7514 2346 7514 4 _025_
rlabel metal2 s 2806 8092 2806 8092 4 _026_
rlabel metal1 s 2438 8840 2438 8840 4 _027_
rlabel metal1 s 4738 9044 4738 9044 4 _028_
rlabel metal1 s 6486 8976 6486 8976 4 _029_
rlabel metal1 s 7084 8942 7084 8942 4 _030_
rlabel metal2 s 8234 8636 8234 8636 4 _031_
rlabel metal2 s 4278 8636 4278 8636 4 _032_
rlabel metal2 s 2530 8636 2530 8636 4 _033_
rlabel metal1 s 2162 8432 2162 8432 4 _034_
rlabel metal1 s 1932 5746 1932 5746 4 _035_
rlabel metal2 s 1886 7684 1886 7684 4 _036_
rlabel metal1 s 2116 8058 2116 8058 4 _037_
rlabel metal1 s 4094 8398 4094 8398 4 _038_
rlabel metal1 s 4186 8330 4186 8330 4 _039_
rlabel metal2 s 5474 8670 5474 8670 4 _040_
rlabel metal1 s 3910 8500 3910 8500 4 _041_
rlabel metal2 s 7590 8058 7590 8058 4 _042_
rlabel metal1 s 6026 8976 6026 8976 4 _043_
rlabel metal1 s 6394 8534 6394 8534 4 _044_
rlabel metal1 s 7176 7922 7176 7922 4 _045_
rlabel metal1 s 6946 7854 6946 7854 4 _046_
rlabel metal2 s 7038 9214 7038 9214 4 _047_
rlabel metal2 s 7222 8330 7222 8330 4 _048_
rlabel metal2 s 7774 8228 7774 8228 4 _049_
rlabel metal2 s 8418 8228 8418 8228 4 _050_
rlabel metal1 s 2116 3978 2116 3978 4 _051_
rlabel metal2 s 2262 5610 2262 5610 4 _052_
rlabel metal2 s 1610 5372 1610 5372 4 _053_
rlabel metal1 s 4554 5202 4554 5202 4 _054_
rlabel metal2 s 4278 5576 4278 5576 4 _055_
rlabel metal1 s 4064 5610 4064 5610 4 _056_
rlabel metal1 s 4094 3944 4094 3944 4 _057_
rlabel metal1 s 4370 4148 4370 4148 4 _058_
rlabel metal2 s 6394 4624 6394 4624 4 _059_
rlabel metal1 s 5750 3910 5750 3910 4 _060_
rlabel metal1 s 5712 4250 5712 4250 4 _061_
rlabel metal2 s 6578 5100 6578 5100 4 _062_
rlabel metal2 s 7866 4318 7866 4318 4 _063_
rlabel metal1 s 7084 4794 7084 4794 4 _064_
rlabel metal1 s 7590 6630 7590 6630 4 _065_
rlabel metal2 s 5842 7140 5842 7140 4 _066_
rlabel metal1 s 3266 7344 3266 7344 4 _067_
rlabel metal1 s 4002 7378 4002 7378 4 _068_
rlabel metal1 s 5566 7344 5566 7344 4 _069_
rlabel metal1 s 5428 6630 5428 6630 4 _070_
rlabel metal2 s 6394 6970 6394 6970 4 _071_
rlabel metal1 s 7314 6766 7314 6766 4 _072_
rlabel metal2 s 4462 5389 4462 5389 4 clk
rlabel metal1 s 4692 5338 4692 5338 4 clknet_0_clk
rlabel metal2 s 1794 4080 1794 4080 4 clknet_1_0__leaf_clk
rlabel metal2 s 6486 3264 6486 3264 4 clknet_1_1__leaf_clk
rlabel metal1 s 1978 6732 1978 6732 4 counter\[0\]
rlabel metal2 s 1794 6562 1794 6562 4 counter\[1\]
rlabel metal2 s 3542 8364 3542 8364 4 counter\[2\]
rlabel metal2 s 4922 6052 4922 6052 4 counter\[3\]
rlabel metal1 s 5428 8466 5428 8466 4 counter\[4\]
rlabel metal1 s 5382 4080 5382 4080 4 counter\[5\]
rlabel metal1 s 7728 4114 7728 4114 4 counter\[6\]
rlabel metal2 s 8602 4828 8602 4828 4 counter\[7\]
rlabel metal1 s 1564 8262 1564 8262 4 net1
rlabel metal2 s 7958 5882 7958 5882 4 net10
rlabel metal1 s 8326 2822 8326 2822 4 net11
rlabel metal1 s 7958 5882 7958 5882 4 net12
rlabel metal1 s 2714 8908 2714 8908 4 net2
rlabel metal1 s 2438 9010 2438 9010 4 net3
rlabel metal2 s 3634 9282 3634 9282 4 net4
rlabel metal1 s 5612 9146 5612 9146 4 net5
rlabel metal2 s 5566 8398 5566 8398 4 net6
rlabel metal2 s 6670 8160 6670 8160 4 net7
rlabel metal1 s 8280 7378 8280 7378 4 net8
rlabel metal2 s 8326 2689 8326 2689 4 net9
rlabel metal1 s 8050 5814 8050 5814 4 out
rlabel metal3 s 1050 8228 1050 8228 4 psc[0]
rlabel metal3 s 0 7488 800 7608 4 psc[1]
port 6 nsew
rlabel metal3 s 0 8848 800 8968 4 psc[2]
port 7 nsew
rlabel metal1 s 4002 9588 4002 9588 4 psc[3]
rlabel metal1 s 5658 9622 5658 9622 4 psc[4]
rlabel metal1 s 5980 9554 5980 9554 4 psc[5]
rlabel metal1 s 6532 9554 6532 9554 4 psc[6]
rlabel metal2 s 8694 7089 8694 7089 4 psc[7]
rlabel metal2 s 8694 3247 8694 3247 4 rst
flabel metal4 s 4868 2128 5188 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4208 2128 4528 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 9405 5448 10205 5568 0 FreeSans 600 0 0 0 out
port 4 nsew
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 psc[0]
port 5 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 psc[1]
flabel metal3 s 400 8908 400 8908 0 FreeSans 600 0 0 0 psc[2]
flabel metal2 s 3238 11549 3294 12349 0 FreeSans 280 90 0 0 psc[3]
port 8 nsew
flabel metal2 s 5170 11549 5226 12349 0 FreeSans 280 90 0 0 psc[4]
port 9 nsew
flabel metal2 s 5814 11549 5870 12349 0 FreeSans 280 90 0 0 psc[5]
port 10 nsew
flabel metal2 s 6458 11549 6514 12349 0 FreeSans 280 90 0 0 psc[6]
port 11 nsew
flabel metal3 s 9405 6808 10205 6928 0 FreeSans 600 0 0 0 psc[7]
port 12 nsew
flabel metal3 s 9405 3408 10205 3528 0 FreeSans 600 0 0 0 rst
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 10205 12349
<< end >>
