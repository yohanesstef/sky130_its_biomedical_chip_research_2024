magic
tech sky130A
magscale 1 2
timestamp 1730527170
<< nmos >>
rect -15 -219 15 281
<< ndiff >>
rect -73 269 -15 281
rect -73 -207 -61 269
rect -27 -207 -15 269
rect -73 -219 -15 -207
rect 15 269 73 281
rect 15 -207 27 269
rect 61 -207 73 269
rect 15 -219 73 -207
<< ndiffc >>
rect -61 -207 -27 269
rect 27 -207 61 269
<< poly >>
rect -15 281 15 307
rect -15 -241 15 -219
rect -33 -257 33 -241
rect -33 -291 -17 -257
rect 17 -291 33 -257
rect -33 -307 33 -291
<< polycont >>
rect -17 -291 17 -257
<< locali >>
rect -61 269 -27 285
rect -61 -223 -27 -207
rect 27 269 61 285
rect 27 -223 61 -207
rect -33 -291 -17 -257
rect 17 -291 33 -257
<< viali >>
rect -61 -207 -27 269
rect 27 -207 61 269
<< metal1 >>
rect -67 269 -21 281
rect -67 -207 -61 269
rect -27 -207 -21 269
rect -67 -219 -21 -207
rect 21 269 67 281
rect 21 -207 27 269
rect 61 -207 67 269
rect 21 -219 67 -207
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
