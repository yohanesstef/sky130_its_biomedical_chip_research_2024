module freq_psc (clk,
    out,
    rst,
    psc);
 input clk;
 output out;
 input rst;
 input [31:0] psc;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire \psc_cnt[0] ;
 wire \psc_cnt[10] ;
 wire \psc_cnt[11] ;
 wire \psc_cnt[12] ;
 wire \psc_cnt[13] ;
 wire \psc_cnt[14] ;
 wire \psc_cnt[15] ;
 wire \psc_cnt[16] ;
 wire \psc_cnt[17] ;
 wire \psc_cnt[18] ;
 wire \psc_cnt[19] ;
 wire \psc_cnt[1] ;
 wire \psc_cnt[20] ;
 wire \psc_cnt[21] ;
 wire \psc_cnt[22] ;
 wire \psc_cnt[23] ;
 wire \psc_cnt[24] ;
 wire \psc_cnt[25] ;
 wire \psc_cnt[26] ;
 wire \psc_cnt[27] ;
 wire \psc_cnt[28] ;
 wire \psc_cnt[29] ;
 wire \psc_cnt[2] ;
 wire \psc_cnt[30] ;
 wire \psc_cnt[31] ;
 wire \psc_cnt[3] ;
 wire \psc_cnt[4] ;
 wire \psc_cnt[5] ;
 wire \psc_cnt[6] ;
 wire \psc_cnt[7] ;
 wire \psc_cnt[8] ;
 wire \psc_cnt[9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net59;

 sky130_fd_sc_hd__inv_2 _236_ (.A(\psc_cnt[24] ),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _237_ (.A(net15),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _238_ (.A(net14),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(\psc_cnt[20] ),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(\psc_cnt[19] ),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(net10),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _242_ (.A(net9),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(net8),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _244_ (.A(\psc_cnt[15] ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _245_ (.A(\psc_cnt[14] ),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(\psc_cnt[13] ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _247_ (.A(\psc_cnt[12] ),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _248_ (.A(\psc_cnt[11] ),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _249_ (.A(\psc_cnt[10] ),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _250_ (.A(\psc_cnt[9] ),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _251_ (.A(\psc_cnt[8] ),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(net31),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(net30),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _254_ (.A(net29),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _255_ (.A(net28),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _256_ (.A(net27),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _257_ (.A(net26),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _258_ (.A(net23),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _259_ (.A(net12),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(net1),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(\psc_cnt[25] ),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _262_ (.A(\psc_cnt[26] ),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(\psc_cnt[28] ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(\psc_cnt[29] ),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _265_ (.A(net43),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(net39),
    .Y(_032_));
 sky130_fd_sc_hd__and2_1 _267_ (.A(net7),
    .B(_074_),
    .X(_096_));
 sky130_fd_sc_hd__o22a_1 _268_ (.A1(net7),
    .A2(_074_),
    .B1(net6),
    .B2(_075_),
    .X(_097_));
 sky130_fd_sc_hd__a22oi_1 _269_ (.A1(net6),
    .A2(_075_),
    .B1(net5),
    .B2(_076_),
    .Y(_098_));
 sky130_fd_sc_hd__o22a_1 _270_ (.A1(net5),
    .A2(_076_),
    .B1(_077_),
    .B2(net4),
    .X(_099_));
 sky130_fd_sc_hd__nand2b_1 _271_ (.A_N(_099_),
    .B(_098_),
    .Y(_100_));
 sky130_fd_sc_hd__a21oi_1 _272_ (.A1(_097_),
    .A2(_100_),
    .B1(_096_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_1 _273_ (.A1(_077_),
    .A2(net4),
    .B1(_096_),
    .Y(_102_));
 sky130_fd_sc_hd__and4_1 _274_ (.A(_097_),
    .B(_098_),
    .C(_099_),
    .D(_102_),
    .X(_103_));
 sky130_fd_sc_hd__and2b_1 _275_ (.A_N(\psc_cnt[11] ),
    .B(net3),
    .X(_104_));
 sky130_fd_sc_hd__o22a_1 _276_ (.A1(net3),
    .A2(_078_),
    .B1(net2),
    .B2(_079_),
    .X(_105_));
 sky130_fd_sc_hd__a221oi_1 _277_ (.A1(net2),
    .A2(_079_),
    .B1(net32),
    .B2(_080_),
    .C1(_104_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_1 _278_ (.A(_105_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__o22a_1 _279_ (.A1(net32),
    .A2(_080_),
    .B1(_081_),
    .B2(net31),
    .X(_108_));
 sky130_fd_sc_hd__a22o_1 _280_ (.A1(_085_),
    .A2(\psc_cnt[5] ),
    .B1(\psc_cnt[4] ),
    .B2(_086_),
    .X(_109_));
 sky130_fd_sc_hd__a211o_1 _281_ (.A1(_089_),
    .A2(\psc_cnt[1] ),
    .B1(_090_),
    .C1(\psc_cnt[0] ),
    .X(_110_));
 sky130_fd_sc_hd__o22a_1 _282_ (.A1(_088_),
    .A2(\psc_cnt[2] ),
    .B1(_089_),
    .B2(\psc_cnt[1] ),
    .X(_111_));
 sky130_fd_sc_hd__a22o_1 _283_ (.A1(_087_),
    .A2(\psc_cnt[3] ),
    .B1(_088_),
    .B2(\psc_cnt[2] ),
    .X(_112_));
 sky130_fd_sc_hd__a21o_1 _284_ (.A1(_110_),
    .A2(_111_),
    .B1(_112_),
    .X(_113_));
 sky130_fd_sc_hd__o22a_1 _285_ (.A1(\psc_cnt[4] ),
    .A2(_086_),
    .B1(_087_),
    .B2(\psc_cnt[3] ),
    .X(_114_));
 sky130_fd_sc_hd__a21o_1 _286_ (.A1(_113_),
    .A2(_114_),
    .B1(_109_),
    .X(_115_));
 sky130_fd_sc_hd__o22a_1 _287_ (.A1(_084_),
    .A2(\psc_cnt[6] ),
    .B1(_085_),
    .B2(\psc_cnt[5] ),
    .X(_116_));
 sky130_fd_sc_hd__a22o_1 _288_ (.A1(_083_),
    .A2(\psc_cnt[7] ),
    .B1(_084_),
    .B2(\psc_cnt[6] ),
    .X(_117_));
 sky130_fd_sc_hd__a21o_1 _289_ (.A1(_115_),
    .A2(_116_),
    .B1(_117_),
    .X(_118_));
 sky130_fd_sc_hd__o221a_1 _290_ (.A1(\psc_cnt[8] ),
    .A2(_082_),
    .B1(_083_),
    .B2(\psc_cnt[7] ),
    .C1(_108_),
    .X(_119_));
 sky130_fd_sc_hd__and4_1 _291_ (.A(_103_),
    .B(_105_),
    .C(_106_),
    .D(_119_),
    .X(_120_));
 sky130_fd_sc_hd__o22a_1 _292_ (.A1(_104_),
    .A2(_105_),
    .B1(_107_),
    .B2(_108_),
    .X(_121_));
 sky130_fd_sc_hd__and2b_1 _293_ (.A_N(_121_),
    .B(_103_),
    .X(_122_));
 sky130_fd_sc_hd__a211o_1 _294_ (.A1(_118_),
    .A2(_120_),
    .B1(_122_),
    .C1(_101_),
    .X(_123_));
 sky130_fd_sc_hd__a2bb2o_1 _295_ (.A1_N(net11),
    .A2_N(_070_),
    .B1(_071_),
    .B2(\psc_cnt[18] ),
    .X(_124_));
 sky130_fd_sc_hd__nand2_1 _296_ (.A(net11),
    .B(_070_),
    .Y(_125_));
 sky130_fd_sc_hd__or2_1 _297_ (.A(_071_),
    .B(\psc_cnt[18] ),
    .X(_126_));
 sky130_fd_sc_hd__and3b_1 _298_ (.A_N(_124_),
    .B(_125_),
    .C(_126_),
    .X(_127_));
 sky130_fd_sc_hd__a22o_1 _299_ (.A1(_072_),
    .A2(\psc_cnt[17] ),
    .B1(\psc_cnt[16] ),
    .B2(_073_),
    .X(_128_));
 sky130_fd_sc_hd__or2_1 _300_ (.A(_072_),
    .B(\psc_cnt[17] ),
    .X(_129_));
 sky130_fd_sc_hd__o21a_1 _301_ (.A1(\psc_cnt[16] ),
    .A2(_073_),
    .B1(_127_),
    .X(_130_));
 sky130_fd_sc_hd__and2b_1 _302_ (.A_N(net16),
    .B(\psc_cnt[23] ),
    .X(_131_));
 sky130_fd_sc_hd__a21o_1 _303_ (.A1(_067_),
    .A2(\psc_cnt[22] ),
    .B1(_131_),
    .X(_132_));
 sky130_fd_sc_hd__and2b_1 _304_ (.A_N(net13),
    .B(\psc_cnt[20] ),
    .X(_133_));
 sky130_fd_sc_hd__and2b_1 _305_ (.A_N(net14),
    .B(\psc_cnt[21] ),
    .X(_134_));
 sky130_fd_sc_hd__a2111o_1 _306_ (.A1(_067_),
    .A2(\psc_cnt[22] ),
    .B1(_131_),
    .C1(_133_),
    .D1(_134_),
    .X(_135_));
 sky130_fd_sc_hd__and2b_1 _307_ (.A_N(net20),
    .B(\psc_cnt[27] ),
    .X(_136_));
 sky130_fd_sc_hd__and2b_1 _308_ (.A_N(net19),
    .B(\psc_cnt[26] ),
    .X(_137_));
 sky130_fd_sc_hd__nor2_1 _309_ (.A(_136_),
    .B(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__and2b_1 _310_ (.A_N(\psc_cnt[27] ),
    .B(net20),
    .X(_139_));
 sky130_fd_sc_hd__and2b_1 _311_ (.A_N(\psc_cnt[26] ),
    .B(net19),
    .X(_140_));
 sky130_fd_sc_hd__or4_1 _312_ (.A(_136_),
    .B(_137_),
    .C(_139_),
    .D(_140_),
    .X(_141_));
 sky130_fd_sc_hd__and2b_1 _313_ (.A_N(\psc_cnt[24] ),
    .B(net17),
    .X(_142_));
 sky130_fd_sc_hd__and2b_1 _314_ (.A_N(\psc_cnt[25] ),
    .B(net18),
    .X(_143_));
 sky130_fd_sc_hd__and2b_1 _315_ (.A_N(\psc_cnt[23] ),
    .B(net16),
    .X(_144_));
 sky130_fd_sc_hd__or3_1 _316_ (.A(_142_),
    .B(_143_),
    .C(_144_),
    .X(_145_));
 sky130_fd_sc_hd__or3_1 _317_ (.A(_135_),
    .B(_141_),
    .C(_145_),
    .X(_146_));
 sky130_fd_sc_hd__and2b_1 _318_ (.A_N(net25),
    .B(\psc_cnt[31] ),
    .X(_147_));
 sky130_fd_sc_hd__and2b_1 _319_ (.A_N(net24),
    .B(\psc_cnt[30] ),
    .X(_148_));
 sky130_fd_sc_hd__nor2_1 _320_ (.A(_147_),
    .B(net45),
    .Y(_149_));
 sky130_fd_sc_hd__and2b_1 _321_ (.A_N(\psc_cnt[31] ),
    .B(net25),
    .X(_150_));
 sky130_fd_sc_hd__and2b_1 _322_ (.A_N(\psc_cnt[30] ),
    .B(net24),
    .X(_151_));
 sky130_fd_sc_hd__and2_1 _323_ (.A(_094_),
    .B(net22),
    .X(_152_));
 sky130_fd_sc_hd__or4_4 _324_ (.A(_151_),
    .B(_148_),
    .C(_150_),
    .D(_147_),
    .X(_153_));
 sky130_fd_sc_hd__nor2_1 _325_ (.A(_152_),
    .B(net47),
    .Y(_154_));
 sky130_fd_sc_hd__o22a_1 _326_ (.A1(_094_),
    .A2(net22),
    .B1(net21),
    .B2(_093_),
    .X(_155_));
 sky130_fd_sc_hd__and2b_1 _327_ (.A_N(\psc_cnt[28] ),
    .B(net21),
    .X(_156_));
 sky130_fd_sc_hd__a21oi_1 _328_ (.A1(_069_),
    .A2(net13),
    .B1(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__o22a_1 _329_ (.A1(_066_),
    .A2(net17),
    .B1(_091_),
    .B2(net18),
    .X(_158_));
 sky130_fd_sc_hd__o22a_1 _330_ (.A1(_067_),
    .A2(\psc_cnt[22] ),
    .B1(_068_),
    .B2(\psc_cnt[21] ),
    .X(_159_));
 sky130_fd_sc_hd__and4_1 _331_ (.A(_155_),
    .B(_157_),
    .C(_158_),
    .D(_159_),
    .X(_160_));
 sky130_fd_sc_hd__or4b_4 _332_ (.A(_152_),
    .B(_156_),
    .C(_153_),
    .D_N(_155_),
    .X(_161_));
 sky130_fd_sc_hd__or4_4 _333_ (.A(_141_),
    .B(_142_),
    .C(_143_),
    .D(_161_),
    .X(_162_));
 sky130_fd_sc_hd__and3b_1 _334_ (.A_N(_146_),
    .B(_154_),
    .C(_160_),
    .X(_163_));
 sky130_fd_sc_hd__and4b_1 _335_ (.A_N(_128_),
    .B(_129_),
    .C(_130_),
    .D(_163_),
    .X(_164_));
 sky130_fd_sc_hd__a32o_1 _336_ (.A1(_127_),
    .A2(_128_),
    .A3(_129_),
    .B1(_125_),
    .B2(_124_),
    .X(_165_));
 sky130_fd_sc_hd__and2_1 _337_ (.A(_163_),
    .B(_165_),
    .X(_166_));
 sky130_fd_sc_hd__o32a_1 _338_ (.A1(_141_),
    .A2(_143_),
    .A3(_158_),
    .B1(_139_),
    .B2(_138_),
    .X(_167_));
 sky130_fd_sc_hd__o32a_1 _339_ (.A1(_152_),
    .A2(net46),
    .A3(_155_),
    .B1(_150_),
    .B2(_149_),
    .X(_168_));
 sky130_fd_sc_hd__o21ai_1 _340_ (.A1(_161_),
    .A2(_167_),
    .B1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__o21ba_1 _341_ (.A1(_132_),
    .A2(_159_),
    .B1_N(_144_),
    .X(_170_));
 sky130_fd_sc_hd__and4b_1 _342_ (.A_N(_162_),
    .B(_135_),
    .C(_158_),
    .D(_170_),
    .X(_171_));
 sky130_fd_sc_hd__or3_4 _343_ (.A(_171_),
    .B(_169_),
    .C(_166_),
    .X(_172_));
 sky130_fd_sc_hd__a21oi_4 _344_ (.A1(_123_),
    .A2(_164_),
    .B1(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__xnor2_1 _345_ (.A(net59),
    .B(net35),
    .Y(_065_));
 sky130_fd_sc_hd__and2b_1 _346_ (.A_N(\psc_cnt[0] ),
    .B(net35),
    .X(_000_));
 sky130_fd_sc_hd__or2_1 _347_ (.A(\psc_cnt[1] ),
    .B(\psc_cnt[0] ),
    .X(_174_));
 sky130_fd_sc_hd__nand2_1 _348_ (.A(\psc_cnt[1] ),
    .B(\psc_cnt[0] ),
    .Y(_175_));
 sky130_fd_sc_hd__and3_1 _349_ (.A(net35),
    .B(_174_),
    .C(_175_),
    .X(_011_));
 sky130_fd_sc_hd__a21o_1 _350_ (.A1(\psc_cnt[1] ),
    .A2(\psc_cnt[0] ),
    .B1(\psc_cnt[2] ),
    .X(_176_));
 sky130_fd_sc_hd__nand3_1 _351_ (.A(\psc_cnt[2] ),
    .B(\psc_cnt[1] ),
    .C(\psc_cnt[0] ),
    .Y(_177_));
 sky130_fd_sc_hd__and3_1 _352_ (.A(net35),
    .B(_176_),
    .C(_177_),
    .X(_022_));
 sky130_fd_sc_hd__a31o_1 _353_ (.A1(\psc_cnt[2] ),
    .A2(\psc_cnt[1] ),
    .A3(\psc_cnt[0] ),
    .B1(\psc_cnt[3] ),
    .X(_178_));
 sky130_fd_sc_hd__and4_1 _354_ (.A(\psc_cnt[3] ),
    .B(\psc_cnt[2] ),
    .C(\psc_cnt[1] ),
    .D(\psc_cnt[0] ),
    .X(_179_));
 sky130_fd_sc_hd__and3b_1 _355_ (.A_N(_179_),
    .B(net36),
    .C(_178_),
    .X(_025_));
 sky130_fd_sc_hd__or2_1 _356_ (.A(\psc_cnt[4] ),
    .B(_179_),
    .X(_180_));
 sky130_fd_sc_hd__nand2_1 _357_ (.A(\psc_cnt[4] ),
    .B(_179_),
    .Y(_181_));
 sky130_fd_sc_hd__and3_1 _358_ (.A(net36),
    .B(_180_),
    .C(_181_),
    .X(_026_));
 sky130_fd_sc_hd__a21o_1 _359_ (.A1(\psc_cnt[4] ),
    .A2(_179_),
    .B1(\psc_cnt[5] ),
    .X(_182_));
 sky130_fd_sc_hd__and2_1 _360_ (.A(\psc_cnt[5] ),
    .B(\psc_cnt[4] ),
    .X(_183_));
 sky130_fd_sc_hd__and2_1 _361_ (.A(_179_),
    .B(_183_),
    .X(_184_));
 sky130_fd_sc_hd__and3b_1 _362_ (.A_N(_184_),
    .B(_182_),
    .C(net38),
    .X(_027_));
 sky130_fd_sc_hd__or2_1 _363_ (.A(\psc_cnt[6] ),
    .B(_184_),
    .X(_185_));
 sky130_fd_sc_hd__nand2_1 _364_ (.A(\psc_cnt[6] ),
    .B(_184_),
    .Y(_186_));
 sky130_fd_sc_hd__and3_1 _365_ (.A(net38),
    .B(_185_),
    .C(_186_),
    .X(_028_));
 sky130_fd_sc_hd__a31o_1 _366_ (.A1(\psc_cnt[6] ),
    .A2(_179_),
    .A3(_183_),
    .B1(\psc_cnt[7] ),
    .X(_187_));
 sky130_fd_sc_hd__and4_1 _367_ (.A(\psc_cnt[7] ),
    .B(\psc_cnt[6] ),
    .C(_179_),
    .D(_183_),
    .X(_188_));
 sky130_fd_sc_hd__and3b_1 _368_ (.A_N(_188_),
    .B(_187_),
    .C(net38),
    .X(_029_));
 sky130_fd_sc_hd__or2_1 _369_ (.A(\psc_cnt[8] ),
    .B(_188_),
    .X(_189_));
 sky130_fd_sc_hd__nand2_1 _370_ (.A(\psc_cnt[8] ),
    .B(_188_),
    .Y(_190_));
 sky130_fd_sc_hd__and3_1 _371_ (.A(net38),
    .B(_189_),
    .C(_190_),
    .X(_030_));
 sky130_fd_sc_hd__nand2_1 _372_ (.A(_080_),
    .B(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__nor2_1 _373_ (.A(_080_),
    .B(_081_),
    .Y(_192_));
 sky130_fd_sc_hd__and2_1 _374_ (.A(_188_),
    .B(_192_),
    .X(_193_));
 sky130_fd_sc_hd__and3b_1 _375_ (.A_N(_193_),
    .B(_191_),
    .C(net38),
    .X(_031_));
 sky130_fd_sc_hd__or2_1 _376_ (.A(\psc_cnt[10] ),
    .B(_193_),
    .X(_194_));
 sky130_fd_sc_hd__and3_1 _377_ (.A(\psc_cnt[10] ),
    .B(_188_),
    .C(_192_),
    .X(_195_));
 sky130_fd_sc_hd__and3b_1 _378_ (.A_N(_195_),
    .B(_194_),
    .C(net38),
    .X(_001_));
 sky130_fd_sc_hd__or2_1 _379_ (.A(\psc_cnt[11] ),
    .B(_195_),
    .X(_196_));
 sky130_fd_sc_hd__and4_1 _380_ (.A(\psc_cnt[11] ),
    .B(\psc_cnt[10] ),
    .C(_188_),
    .D(_192_),
    .X(_197_));
 sky130_fd_sc_hd__and3b_1 _381_ (.A_N(_197_),
    .B(net38),
    .C(_196_),
    .X(_002_));
 sky130_fd_sc_hd__and2_1 _382_ (.A(\psc_cnt[12] ),
    .B(_197_),
    .X(_198_));
 sky130_fd_sc_hd__or2_1 _383_ (.A(\psc_cnt[12] ),
    .B(_197_),
    .X(_199_));
 sky130_fd_sc_hd__and3b_1 _384_ (.A_N(_198_),
    .B(_199_),
    .C(net38),
    .X(_003_));
 sky130_fd_sc_hd__or2_1 _385_ (.A(\psc_cnt[13] ),
    .B(_198_),
    .X(_200_));
 sky130_fd_sc_hd__and3_1 _386_ (.A(\psc_cnt[13] ),
    .B(\psc_cnt[12] ),
    .C(_197_),
    .X(_201_));
 sky130_fd_sc_hd__and3b_1 _387_ (.A_N(_201_),
    .B(net37),
    .C(_200_),
    .X(_004_));
 sky130_fd_sc_hd__or2_1 _388_ (.A(\psc_cnt[14] ),
    .B(_201_),
    .X(_202_));
 sky130_fd_sc_hd__nand2_1 _389_ (.A(\psc_cnt[14] ),
    .B(_201_),
    .Y(_203_));
 sky130_fd_sc_hd__and3_1 _390_ (.A(net44),
    .B(_202_),
    .C(_203_),
    .X(_005_));
 sky130_fd_sc_hd__nor2_1 _391_ (.A(_074_),
    .B(_075_),
    .Y(_204_));
 sky130_fd_sc_hd__and4_2 _392_ (.A(\psc_cnt[13] ),
    .B(\psc_cnt[12] ),
    .C(_197_),
    .D(_204_),
    .X(_205_));
 sky130_fd_sc_hd__nand2_1 _393_ (.A(_074_),
    .B(_203_),
    .Y(_206_));
 sky130_fd_sc_hd__and3b_1 _394_ (.A_N(_205_),
    .B(net37),
    .C(_206_),
    .X(_006_));
 sky130_fd_sc_hd__or2_1 _395_ (.A(\psc_cnt[16] ),
    .B(_205_),
    .X(_207_));
 sky130_fd_sc_hd__and2_1 _396_ (.A(\psc_cnt[16] ),
    .B(_205_),
    .X(_208_));
 sky130_fd_sc_hd__and3b_1 _397_ (.A_N(_208_),
    .B(net36),
    .C(_207_),
    .X(_007_));
 sky130_fd_sc_hd__and3_1 _398_ (.A(\psc_cnt[17] ),
    .B(\psc_cnt[16] ),
    .C(_205_),
    .X(_209_));
 sky130_fd_sc_hd__or2_1 _399_ (.A(\psc_cnt[17] ),
    .B(_208_),
    .X(_210_));
 sky130_fd_sc_hd__and3b_1 _400_ (.A_N(_209_),
    .B(_210_),
    .C(net36),
    .X(_008_));
 sky130_fd_sc_hd__nand2_1 _401_ (.A(\psc_cnt[18] ),
    .B(_209_),
    .Y(_211_));
 sky130_fd_sc_hd__o211a_1 _402_ (.A1(\psc_cnt[18] ),
    .A2(_209_),
    .B1(_211_),
    .C1(net36),
    .X(_009_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(_070_),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__and4_1 _404_ (.A(\psc_cnt[19] ),
    .B(\psc_cnt[18] ),
    .C(\psc_cnt[17] ),
    .D(\psc_cnt[16] ),
    .X(_213_));
 sky130_fd_sc_hd__and2_1 _405_ (.A(_205_),
    .B(_213_),
    .X(_214_));
 sky130_fd_sc_hd__and3b_1 _406_ (.A_N(_214_),
    .B(net35),
    .C(_212_),
    .X(_010_));
 sky130_fd_sc_hd__or2_1 _407_ (.A(\psc_cnt[20] ),
    .B(_214_),
    .X(_215_));
 sky130_fd_sc_hd__and3_1 _408_ (.A(\psc_cnt[20] ),
    .B(_205_),
    .C(_213_),
    .X(_216_));
 sky130_fd_sc_hd__and3b_1 _409_ (.A_N(_216_),
    .B(net35),
    .C(_215_),
    .X(_012_));
 sky130_fd_sc_hd__nand2_1 _410_ (.A(\psc_cnt[21] ),
    .B(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__o211a_1 _411_ (.A1(\psc_cnt[21] ),
    .A2(_216_),
    .B1(_217_),
    .C1(net35),
    .X(_013_));
 sky130_fd_sc_hd__a21o_1 _412_ (.A1(\psc_cnt[21] ),
    .A2(_216_),
    .B1(\psc_cnt[22] ),
    .X(_218_));
 sky130_fd_sc_hd__and3_1 _413_ (.A(\psc_cnt[22] ),
    .B(\psc_cnt[21] ),
    .C(\psc_cnt[20] ),
    .X(_219_));
 sky130_fd_sc_hd__nand2_1 _414_ (.A(_214_),
    .B(_219_),
    .Y(_220_));
 sky130_fd_sc_hd__and3_1 _415_ (.A(net35),
    .B(_218_),
    .C(_220_),
    .X(_014_));
 sky130_fd_sc_hd__a31o_1 _416_ (.A1(_205_),
    .A2(_213_),
    .A3(_219_),
    .B1(\psc_cnt[23] ),
    .X(_221_));
 sky130_fd_sc_hd__and3_1 _417_ (.A(\psc_cnt[23] ),
    .B(_213_),
    .C(_219_),
    .X(_222_));
 sky130_fd_sc_hd__and2_1 _418_ (.A(_205_),
    .B(_222_),
    .X(_223_));
 sky130_fd_sc_hd__and3b_1 _419_ (.A_N(_223_),
    .B(net35),
    .C(_221_),
    .X(_015_));
 sky130_fd_sc_hd__or2_1 _420_ (.A(\psc_cnt[24] ),
    .B(_223_),
    .X(_224_));
 sky130_fd_sc_hd__and3_1 _421_ (.A(\psc_cnt[24] ),
    .B(_205_),
    .C(_222_),
    .X(_225_));
 sky130_fd_sc_hd__and3b_1 _422_ (.A_N(_225_),
    .B(net35),
    .C(_224_),
    .X(_016_));
 sky130_fd_sc_hd__nand2_1 _423_ (.A(\psc_cnt[25] ),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__o211a_1 _424_ (.A1(\psc_cnt[25] ),
    .A2(_225_),
    .B1(_226_),
    .C1(net44),
    .X(_017_));
 sky130_fd_sc_hd__nand2_1 _425_ (.A(_092_),
    .B(_226_),
    .Y(_227_));
 sky130_fd_sc_hd__o211a_1 _426_ (.A1(_092_),
    .A2(_226_),
    .B1(_227_),
    .C1(net44),
    .X(_018_));
 sky130_fd_sc_hd__a31o_1 _427_ (.A1(\psc_cnt[25] ),
    .A2(\psc_cnt[26] ),
    .A3(_225_),
    .B1(\psc_cnt[27] ),
    .X(_228_));
 sky130_fd_sc_hd__and4_1 _428_ (.A(\psc_cnt[24] ),
    .B(\psc_cnt[25] ),
    .C(\psc_cnt[26] ),
    .D(\psc_cnt[27] ),
    .X(_229_));
 sky130_fd_sc_hd__and3_1 _429_ (.A(_205_),
    .B(_222_),
    .C(_229_),
    .X(_230_));
 sky130_fd_sc_hd__and3b_1 _430_ (.A_N(_230_),
    .B(net37),
    .C(_228_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_1 _431_ (.A(\psc_cnt[28] ),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__o211a_1 _432_ (.A1(\psc_cnt[28] ),
    .A2(_230_),
    .B1(_231_),
    .C1(net44),
    .X(_020_));
 sky130_fd_sc_hd__nand2_1 _433_ (.A(_094_),
    .B(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__and3_1 _434_ (.A(\psc_cnt[28] ),
    .B(\psc_cnt[29] ),
    .C(_230_),
    .X(_233_));
 sky130_fd_sc_hd__and3b_1 _435_ (.A_N(_233_),
    .B(net37),
    .C(_232_),
    .X(_021_));
 sky130_fd_sc_hd__or2_1 _436_ (.A(\psc_cnt[30] ),
    .B(_233_),
    .X(_234_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(\psc_cnt[30] ),
    .B(_233_),
    .Y(_235_));
 sky130_fd_sc_hd__and3_1 _438_ (.A(net37),
    .B(_234_),
    .C(_235_),
    .X(_023_));
 sky130_fd_sc_hd__a21boi_1 _439_ (.A1(_095_),
    .A2(_235_),
    .B1_N(net44),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _440_ (.A(net39),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _441_ (.A(net40),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _442_ (.A(net40),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _443_ (.A(net40),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _444_ (.A(net41),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _445_ (.A(net42),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _446_ (.A(net42),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _447_ (.A(net42),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _448_ (.A(net42),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _449_ (.A(net42),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _450_ (.A(net42),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _451_ (.A(net42),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _452_ (.A(net41),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _453_ (.A(net41),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _454_ (.A(net41),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _455_ (.A(net40),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _456_ (.A(net40),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _457_ (.A(net40),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _458_ (.A(net39),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _459_ (.A(net39),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _460_ (.A(net39),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _461_ (.A(net39),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _462_ (.A(net39),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _463_ (.A(net39),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _464_ (.A(net39),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _465_ (.A(net41),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _466_ (.A(net41),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _467_ (.A(net41),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _468_ (.A(net41),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _469_ (.A(net41),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _470_ (.A(net41),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _471_ (.A(net39),
    .Y(_064_));
 sky130_fd_sc_hd__dfrtp_2 _472_ (.CLK(clknet_2_1__leaf_clk),
    .D(_000_),
    .RESET_B(_032_),
    .Q(\psc_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _473_ (.CLK(clknet_2_1__leaf_clk),
    .D(_011_),
    .RESET_B(_033_),
    .Q(\psc_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _474_ (.CLK(clknet_2_1__leaf_clk),
    .D(_022_),
    .RESET_B(_034_),
    .Q(\psc_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _475_ (.CLK(clknet_2_1__leaf_clk),
    .D(_025_),
    .RESET_B(_035_),
    .Q(\psc_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _476_ (.CLK(clknet_2_1__leaf_clk),
    .D(_026_),
    .RESET_B(_036_),
    .Q(\psc_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _477_ (.CLK(clknet_2_1__leaf_clk),
    .D(_027_),
    .RESET_B(_037_),
    .Q(\psc_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _478_ (.CLK(clknet_2_3__leaf_clk),
    .D(_028_),
    .RESET_B(_038_),
    .Q(\psc_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _479_ (.CLK(clknet_2_3__leaf_clk),
    .D(_029_),
    .RESET_B(_039_),
    .Q(\psc_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _480_ (.CLK(clknet_2_3__leaf_clk),
    .D(_030_),
    .RESET_B(_040_),
    .Q(\psc_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _481_ (.CLK(clknet_2_3__leaf_clk),
    .D(_031_),
    .RESET_B(_041_),
    .Q(\psc_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _482_ (.CLK(clknet_2_3__leaf_clk),
    .D(_001_),
    .RESET_B(_042_),
    .Q(\psc_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _483_ (.CLK(clknet_2_3__leaf_clk),
    .D(_002_),
    .RESET_B(_043_),
    .Q(\psc_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _484_ (.CLK(clknet_2_3__leaf_clk),
    .D(_003_),
    .RESET_B(_044_),
    .Q(\psc_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _485_ (.CLK(clknet_2_2__leaf_clk),
    .D(_004_),
    .RESET_B(_045_),
    .Q(\psc_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _486_ (.CLK(clknet_2_2__leaf_clk),
    .D(_005_),
    .RESET_B(_046_),
    .Q(\psc_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _487_ (.CLK(clknet_2_2__leaf_clk),
    .D(_006_),
    .RESET_B(_047_),
    .Q(\psc_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _488_ (.CLK(clknet_2_1__leaf_clk),
    .D(_007_),
    .RESET_B(_048_),
    .Q(\psc_cnt[16] ));
 sky130_fd_sc_hd__dfrtp_1 _489_ (.CLK(clknet_2_1__leaf_clk),
    .D(_008_),
    .RESET_B(_049_),
    .Q(\psc_cnt[17] ));
 sky130_fd_sc_hd__dfrtp_1 _490_ (.CLK(clknet_2_0__leaf_clk),
    .D(_009_),
    .RESET_B(_050_),
    .Q(\psc_cnt[18] ));
 sky130_fd_sc_hd__dfrtp_1 _491_ (.CLK(clknet_2_0__leaf_clk),
    .D(_010_),
    .RESET_B(_051_),
    .Q(\psc_cnt[19] ));
 sky130_fd_sc_hd__dfrtp_1 _492_ (.CLK(clknet_2_0__leaf_clk),
    .D(_012_),
    .RESET_B(_052_),
    .Q(\psc_cnt[20] ));
 sky130_fd_sc_hd__dfrtp_1 _493_ (.CLK(clknet_2_0__leaf_clk),
    .D(_013_),
    .RESET_B(_053_),
    .Q(\psc_cnt[21] ));
 sky130_fd_sc_hd__dfrtp_1 _494_ (.CLK(clknet_2_0__leaf_clk),
    .D(_014_),
    .RESET_B(_054_),
    .Q(\psc_cnt[22] ));
 sky130_fd_sc_hd__dfrtp_1 _495_ (.CLK(clknet_2_0__leaf_clk),
    .D(_015_),
    .RESET_B(_055_),
    .Q(\psc_cnt[23] ));
 sky130_fd_sc_hd__dfrtp_1 _496_ (.CLK(clknet_2_1__leaf_clk),
    .D(_016_),
    .RESET_B(_056_),
    .Q(\psc_cnt[24] ));
 sky130_fd_sc_hd__dfrtp_2 _497_ (.CLK(clknet_2_2__leaf_clk),
    .D(_017_),
    .RESET_B(_057_),
    .Q(\psc_cnt[25] ));
 sky130_fd_sc_hd__dfrtp_1 _498_ (.CLK(clknet_2_2__leaf_clk),
    .D(_018_),
    .RESET_B(_058_),
    .Q(\psc_cnt[26] ));
 sky130_fd_sc_hd__dfrtp_1 _499_ (.CLK(clknet_2_2__leaf_clk),
    .D(_019_),
    .RESET_B(_059_),
    .Q(\psc_cnt[27] ));
 sky130_fd_sc_hd__dfrtp_1 _500_ (.CLK(clknet_2_2__leaf_clk),
    .D(_020_),
    .RESET_B(_060_),
    .Q(\psc_cnt[28] ));
 sky130_fd_sc_hd__dfrtp_1 _501_ (.CLK(clknet_2_2__leaf_clk),
    .D(_021_),
    .RESET_B(_061_),
    .Q(\psc_cnt[29] ));
 sky130_fd_sc_hd__dfrtp_1 _502_ (.CLK(clknet_2_2__leaf_clk),
    .D(_023_),
    .RESET_B(_062_),
    .Q(\psc_cnt[30] ));
 sky130_fd_sc_hd__dfrtp_1 _503_ (.CLK(clknet_2_2__leaf_clk),
    .D(_024_),
    .RESET_B(_063_),
    .Q(\psc_cnt[31] ));
 sky130_fd_sc_hd__dfrtp_1 _504_ (.CLK(clknet_2_0__leaf_clk),
    .D(_065_),
    .RESET_B(_064_),
    .Q(net34));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_121 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(psc[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(psc[10]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(psc[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(psc[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(psc[13]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(psc[14]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(psc[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(psc[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(psc[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(psc[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(psc[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(psc[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(psc[20]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(psc[21]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(psc[22]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(psc[23]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(psc[24]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(psc[25]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(psc[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(psc[27]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(psc[28]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(psc[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(psc[2]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(psc[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(psc[31]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(psc[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(psc[4]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(psc[5]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(psc[6]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(psc[7]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(psc[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(psc[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(rst),
    .X(net33));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(out));
 sky130_fd_sc_hd__buf_6 fanout35 (.A(_173_),
    .X(net35));
 sky130_fd_sc_hd__buf_6 fanout36 (.A(_173_),
    .X(net36));
 sky130_fd_sc_hd__buf_6 fanout37 (.A(_173_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(_173_),
    .X(net38));
 sky130_fd_sc_hd__buf_4 fanout39 (.A(net33),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net33),
    .X(net40));
 sky130_fd_sc_hd__buf_4 fanout41 (.A(net33),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net33),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload0 (.A(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload2 (.A(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(\psc_cnt[31] ),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 clone2 (.A(_173_),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer3 (.A(_148_),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer4 (.A(_153_),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(_153_),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net34),
    .X(net59));
endmodule
