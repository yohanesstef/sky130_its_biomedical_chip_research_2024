magic
tech sky130A
magscale 1 2
timestamp 1729853601
<< error_p >>
rect -32 137 32 143
rect -32 103 -20 137
rect -32 97 32 103
<< pwell >>
rect -232 -275 232 275
<< nmos >>
rect -36 -127 36 65
<< ndiff >>
rect -94 53 -36 65
rect -94 -115 -82 53
rect -48 -115 -36 53
rect -94 -127 -36 -115
rect 36 53 94 65
rect 36 -115 48 53
rect 82 -115 94 53
rect 36 -127 94 -115
<< ndiffc >>
rect -82 -115 -48 53
rect 48 -115 82 53
<< psubdiff >>
rect -196 205 -100 239
rect 100 205 196 239
rect -196 143 -162 205
rect 162 143 196 205
rect -196 -205 -162 -143
rect 162 -205 196 -143
rect -196 -239 -100 -205
rect 100 -239 196 -205
<< psubdiffcont >>
rect -100 205 100 239
rect -196 -143 -162 143
rect 162 -143 196 143
rect -100 -239 100 -205
<< poly >>
rect -36 137 36 153
rect -36 103 -20 137
rect 20 103 36 137
rect -36 65 36 103
rect -36 -153 36 -127
<< polycont >>
rect -20 103 20 137
<< locali >>
rect -196 205 -100 239
rect 100 205 196 239
rect -196 143 -162 205
rect 162 143 196 205
rect -36 103 -20 137
rect 20 103 36 137
rect -82 53 -48 69
rect -82 -131 -48 -115
rect 48 53 82 69
rect 48 -131 82 -115
rect -196 -205 -162 -143
rect 162 -205 196 -143
rect -196 -239 -100 -205
rect 100 -239 196 -205
<< viali >>
rect -20 103 20 137
rect -82 -115 -48 53
rect 48 -115 82 53
<< metal1 >>
rect -32 137 32 143
rect -32 103 -20 137
rect 20 103 32 137
rect -32 97 32 103
rect -88 53 -42 65
rect -88 -115 -82 53
rect -48 -115 -42 53
rect -88 -127 -42 -115
rect 42 53 88 65
rect 42 -115 48 53
rect 82 -115 88 53
rect 42 -127 88 -115
<< properties >>
string FIXED_BBOX -179 -222 179 222
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.96 l 0.36 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
