magic
tech sky130A
timestamp 1729851530
<< nwell >>
rect -56 -271 56 271
<< pmos >>
rect -9 -240 9 240
<< pdiff >>
rect -38 234 -9 240
rect -38 -234 -32 234
rect -15 -234 -9 234
rect -38 -240 -9 -234
rect 9 234 38 240
rect 9 -234 15 234
rect 32 -234 38 234
rect 9 -240 38 -234
<< pdiffc >>
rect -32 -234 -15 234
rect 15 -234 32 234
<< poly >>
rect -9 240 9 253
rect -9 -253 9 -240
<< locali >>
rect -32 234 -15 242
rect -32 -242 -15 -234
rect 15 234 32 242
rect 15 -242 32 -234
<< viali >>
rect -32 -234 -15 234
rect 15 -234 32 234
<< metal1 >>
rect -35 234 -12 240
rect -35 -234 -32 234
rect -15 -234 -12 234
rect -35 -240 -12 -234
rect 12 234 35 240
rect 12 -234 15 234
rect 32 -234 35 234
rect 12 -240 35 -234
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.8 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
