magic
tech sky130A
magscale 1 2
timestamp 1730019635
<< error_p >>
rect -29 -137 29 -131
rect -29 -171 -17 -137
rect -29 -177 29 -171
<< nwell >>
rect -109 -190 109 224
<< pmos >>
rect -15 -90 15 162
<< pdiff >>
rect -73 150 -15 162
rect -73 -78 -61 150
rect -27 -78 -15 150
rect -73 -90 -15 -78
rect 15 150 73 162
rect 15 -78 27 150
rect 61 -78 73 150
rect 15 -90 73 -78
<< pdiffc >>
rect -61 -78 -27 150
rect 27 -78 61 150
<< poly >>
rect -15 162 15 188
rect -15 -121 15 -90
rect -33 -137 33 -121
rect -33 -171 -17 -137
rect 17 -171 33 -137
rect -33 -187 33 -171
<< polycont >>
rect -17 -171 17 -137
<< locali >>
rect -61 150 -27 166
rect -61 -94 -27 -78
rect 27 150 61 166
rect 27 -94 61 -78
rect -33 -171 -17 -137
rect 17 -171 33 -137
<< viali >>
rect -61 -78 -27 150
rect 27 -78 61 150
rect -17 -171 17 -137
<< metal1 >>
rect -67 150 -21 162
rect -67 -78 -61 150
rect -27 -78 -21 150
rect -67 -90 -21 -78
rect 21 150 67 162
rect 21 -78 27 150
rect 61 -78 67 150
rect 21 -90 67 -78
rect -29 -137 29 -131
rect -29 -171 -17 -137
rect 17 -171 29 -137
rect -29 -177 29 -171
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
