magic
tech sky130A
magscale 1 2
timestamp 1730127321
<< nwell >>
rect -214 -1100 214 1100
<< pmos >>
rect -120 -1000 120 1000
<< pdiff >>
rect -178 988 -120 1000
rect -178 -988 -166 988
rect -132 -988 -120 988
rect -178 -1000 -120 -988
rect 120 988 178 1000
rect 120 -988 132 988
rect 166 -988 178 988
rect 120 -1000 178 -988
<< pdiffc >>
rect -166 -988 -132 988
rect 132 -988 166 988
<< poly >>
rect -120 1081 120 1097
rect -120 1047 -104 1081
rect 104 1047 120 1081
rect -120 1000 120 1047
rect -120 -1047 120 -1000
rect -120 -1081 -104 -1047
rect 104 -1081 120 -1047
rect -120 -1097 120 -1081
<< polycont >>
rect -104 1047 104 1081
rect -104 -1081 104 -1047
<< locali >>
rect -120 1047 -104 1081
rect 104 1047 120 1081
rect -166 988 -132 1004
rect -166 -1004 -132 -988
rect 132 988 166 1004
rect 132 -1004 166 -988
rect -120 -1081 -104 -1047
rect 104 -1081 120 -1047
<< viali >>
rect -104 1047 104 1081
rect -166 -988 -132 988
rect 132 -988 166 988
rect -104 -1081 104 -1047
<< metal1 >>
rect -116 1081 116 1087
rect -116 1047 -104 1081
rect 104 1047 116 1081
rect -116 1041 116 1047
rect -172 988 -126 1000
rect -172 -988 -166 988
rect -132 -988 -126 988
rect -172 -1000 -126 -988
rect 126 988 172 1000
rect 126 -988 132 988
rect 166 -988 172 988
rect 126 -1000 172 -988
rect -116 -1047 116 -1041
rect -116 -1081 -104 -1047
rect 104 -1081 116 -1047
rect -116 -1087 116 -1081
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
