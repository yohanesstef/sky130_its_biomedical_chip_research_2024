magic
tech sky130A
timestamp 1730525663
<< nmos >>
rect -60 -125 60 125
<< ndiff >>
rect -89 119 -60 125
rect -89 -119 -83 119
rect -66 -119 -60 119
rect -89 -125 -60 -119
rect 60 119 89 125
rect 60 -119 66 119
rect 83 -119 89 119
rect 60 -125 89 -119
<< ndiffc >>
rect -83 -119 -66 119
rect 66 -119 83 119
<< poly >>
rect -60 161 60 169
rect -60 144 -52 161
rect 52 144 60 161
rect -60 125 60 144
rect -60 -144 60 -125
rect -60 -161 -52 -144
rect 52 -161 60 -144
rect -60 -169 60 -161
<< polycont >>
rect -52 144 52 161
rect -52 -161 52 -144
<< locali >>
rect -60 144 -52 161
rect 52 144 60 161
rect -83 119 -66 127
rect -83 -127 -66 -119
rect 66 119 83 127
rect 66 -127 83 -119
rect -60 -161 -52 -144
rect 52 -161 60 -144
<< viali >>
rect -26 144 26 161
rect -83 -119 -66 119
rect 66 -119 83 119
rect -26 -161 26 -144
<< metal1 >>
rect -32 161 32 164
rect -32 144 -26 161
rect 26 144 32 161
rect -32 141 32 144
rect -86 119 -63 125
rect -86 -119 -83 119
rect -66 -119 -63 119
rect -86 -125 -63 -119
rect 63 119 86 125
rect 63 -119 66 119
rect 83 -119 86 119
rect 63 -125 86 -119
rect -32 -144 32 -141
rect -32 -161 -26 -144
rect 26 -161 32 -144
rect -32 -164 32 -161
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2.5 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
