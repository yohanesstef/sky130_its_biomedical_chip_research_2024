* NGSPICE file created from freq_psc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

.subckt freq_psc VGND VPWR clk out psc[0] psc[10] psc[11] psc[12] psc[13] psc[14]
+ psc[15] psc[16] psc[17] psc[18] psc[19] psc[1] psc[20] psc[21] psc[22] psc[23] psc[24]
+ psc[25] psc[26] psc[27] psc[28] psc[29] psc[2] psc[30] psc[31] psc[3] psc[4] psc[5]
+ psc[6] psc[7] psc[8] psc[9] rst
XTAP_TAPCELL_ROW_24_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_432_ _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__inv_2
XFILLER_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_501_ net6 _103_ _104_ net7 VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__o31a_1
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_415_ net42 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
XFILLER_2_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_680_ _087_ counter\[17\] VGND VGND VPWR VPWR _327_ sky130_fd_sc_hd__and2_1
X_663_ _305_ _306_ _308_ _309_ VGND VGND VPWR VPWR _310_ sky130_fd_sc_hd__and4bb_1
X_732_ _091_ counter\[30\] _306_ _308_ VGND VGND VPWR VPWR _379_ sky130_fd_sc_hd__o22ai_1
X_801_ clknet_2_3__leaf_clk _020_ _062_ VGND VGND VPWR VPWR counter\[28\] sky130_fd_sc_hd__dfrtp_1
X_594_ counter\[10\] _261_ VGND VGND VPWR VPWR _263_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_16_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_646_ counter\[27\] _295_ VGND VGND VPWR VPWR _298_ sky130_fd_sc_hd__nand2_1
X_577_ counter\[5\] counter\[4\] _247_ VGND VGND VPWR VPWR _251_ sky130_fd_sc_hd__and3_1
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_715_ counter\[15\] _089_ VGND VGND VPWR VPWR _362_ sky130_fd_sc_hd__nor2_1
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_431_ net15 net14 _108_ _109_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__or4_2
XFILLER_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_500_ _171_ _178_ VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__nor2_1
X_629_ net36 _285_ _286_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_19_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_414_ counter\[26\] VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__inv_2
XFILLER_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_662_ _091_ counter\[30\] _093_ net21 _307_ VGND VGND VPWR VPWR _309_ sky130_fd_sc_hd__o221a_1
X_800_ clknet_2_3__leaf_clk _019_ _061_ VGND VGND VPWR VPWR counter\[27\] sky130_fd_sc_hd__dfrtp_2
X_731_ _313_ _314_ _311_ VGND VGND VPWR VPWR _378_ sky130_fd_sc_hd__o21bai_1
X_593_ counter\[7\] counter\[10\] _253_ _260_ VGND VGND VPWR VPWR _262_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_27_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_645_ counter\[27\] _295_ VGND VGND VPWR VPWR _297_ sky130_fd_sc_hd__or2_1
X_576_ net54 _249_ _250_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and3_1
X_714_ net4 counter\[11\] VGND VGND VPWR VPWR _361_ sky130_fd_sc_hd__and2b_1
X_430_ net10 net9 VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__or2_1
X_628_ counter\[21\] _283_ VGND VGND VPWR VPWR _286_ sky130_fd_sc_hd__nand2_1
X_559_ counter\[19\] _167_ _169_ counter\[18\] _225_ VGND VGND VPWR VPWR _238_ sky130_fd_sc_hd__a221o_1
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_413_ counter\[27\] VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_20_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_661_ _090_ counter\[29\] counter\[28\] _078_ VGND VGND VPWR VPWR _308_ sky130_fd_sc_hd__o22a_1
X_730_ _332_ _376_ _316_ VGND VGND VPWR VPWR _377_ sky130_fd_sc_hd__o21a_1
X_592_ _261_ net35 _259_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and3b_1
XFILLER_19_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xrebuffer19 counter\[8\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd1_1
X_644_ _295_ _296_ net38 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__and3b_1
X_575_ counter\[4\] _247_ VGND VGND VPWR VPWR _250_ sky130_fd_sc_hd__or2_1
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_713_ net3 _076_ _077_ net2 _359_ VGND VGND VPWR VPWR _360_ sky130_fd_sc_hd__o221a_1
XFILLER_31_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_627_ counter\[21\] _283_ VGND VGND VPWR VPWR _285_ sky130_fd_sc_hd__or2_1
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_558_ _224_ _233_ _234_ _236_ VGND VGND VPWR VPWR _237_ sky130_fd_sc_hd__a31oi_1
X_489_ net9 net8 _107_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__or3_4
X_412_ counter\[30\] VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_660_ _091_ counter\[30\] counter\[31\] VGND VGND VPWR VPWR _307_ sky130_fd_sc_hd__a21oi_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_591_ counter\[7\] _253_ _260_ VGND VGND VPWR VPWR _261_ sky130_fd_sc_hd__and3_1
XFILLER_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_789_ clknet_2_1__leaf_clk _007_ _050_ VGND VGND VPWR VPWR counter\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput34 net34 VGND VGND VPWR VPWR out sky130_fd_sc_hd__buf_2
X_712_ counter\[11\] net4 VGND VGND VPWR VPWR _359_ sky130_fd_sc_hd__nand2b_1
X_574_ counter\[4\] _247_ VGND VGND VPWR VPWR _249_ sky130_fd_sc_hd__nand2_1
X_643_ counter\[26\] _294_ VGND VGND VPWR VPWR _296_ sky130_fd_sc_hd__or2_1
XFILLER_30_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_557_ counter\[15\] _181_ _235_ VGND VGND VPWR VPWR _236_ sky130_fd_sc_hd__o21a_1
X_488_ net11 _152_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__xnor2_2
X_626_ _283_ _284_ net36 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and3b_1
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_411_ net25 VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_609_ counter\[15\] counter\[14\] _269_ VGND VGND VPWR VPWR _273_ sky130_fd_sc_hd__and3_1
XFILLER_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload0 clknet_2_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__bufinv_16
X_590_ counter\[9\] counter\[8\] VGND VGND VPWR VPWR _260_ sky130_fd_sc_hd__and2_1
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_788_ clknet_2_1__leaf_clk _006_ _049_ VGND VGND VPWR VPWR counter\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_573_ _247_ _248_ net37 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and3b_1
X_642_ counter\[26\] counter\[25\] counter\[24\] _290_ VGND VGND VPWR VPWR _295_ sky130_fd_sc_hd__and4_1
XFILLER_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_711_ net5 _075_ VGND VGND VPWR VPWR _358_ sky130_fd_sc_hd__and2_1
XFILLER_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_625_ counter\[20\] _282_ VGND VGND VPWR VPWR _284_ sky130_fd_sc_hd__or2_1
X_487_ counter\[20\] _164_ _165_ VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_14_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_556_ _186_ _189_ _183_ VGND VGND VPWR VPWR _235_ sky130_fd_sc_hd__a21o_1
XFILLER_8_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_410_ net24 VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__inv_2
X_608_ counter\[14\] _269_ counter\[15\] VGND VGND VPWR VPWR _272_ sky130_fd_sc_hd__a21o_1
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_539_ counter\[11\] _191_ _192_ counter\[10\] VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__o22a_1
XFILLER_23_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_2_1__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_29_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_787_ clknet_2_1__leaf_clk _005_ _048_ VGND VGND VPWR VPWR counter\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_25_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_572_ counter\[3\] _245_ VGND VGND VPWR VPWR _248_ sky130_fd_sc_hd__or2_1
X_641_ _294_ net38 _293_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__and3b_1
X_710_ _356_ VGND VGND VPWR VPWR _357_ sky130_fd_sc_hd__inv_2
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_486_ counter\[21\] _160_ _164_ counter\[20\] VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__a22oi_1
X_555_ counter\[15\] _181_ _188_ counter\[12\] _186_ VGND VGND VPWR VPWR _234_ sky130_fd_sc_hd__o221a_1
XFILLER_8_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_624_ counter\[20\] counter\[19\] counter\[18\] _277_ VGND VGND VPWR VPWR _283_ sky130_fd_sc_hd__and4_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_538_ counter\[7\] _198_ _214_ counter\[6\] VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__a22o_1
X_607_ net35 _270_ _271_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__and3_1
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_469_ counter\[27\] _116_ _140_ VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__and3_1
XFILLER_13_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload2 clknet_2_2__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_18_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_786_ clknet_2_0__leaf_clk _004_ _047_ VGND VGND VPWR VPWR counter\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_571_ counter\[0\] counter\[1\] counter\[3\] counter\[2\] VGND VGND VPWR VPWR _247_
+ sky130_fd_sc_hd__and4_1
X_640_ counter\[25\] counter\[24\] _290_ VGND VGND VPWR VPWR _294_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_769_ net43 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__inv_2
XFILLER_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_485_ _153_ _163_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__nor2_1
XFILLER_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_554_ _183_ _189_ VGND VGND VPWR VPWR _233_ sky130_fd_sc_hd__nor2_1
X_623_ _282_ net36 _281_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_20_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_468_ _141_ _143_ _144_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__and3_1
X_399_ net21 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__inv_2
X_537_ counter\[5\] _211_ _212_ _210_ _215_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__o221a_1
X_606_ counter\[14\] _269_ VGND VGND VPWR VPWR _271_ sky130_fd_sc_hd__or2_1
XFILLER_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_785_ clknet_2_0__leaf_clk _003_ _046_ VGND VGND VPWR VPWR counter\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_570_ _245_ _246_ net37 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__and3b_1
XFILLER_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_699_ _067_ net23 VGND VGND VPWR VPWR _346_ sky130_fd_sc_hd__nand2_1
X_768_ net43 VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__inv_2
XFILLER_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_553_ _148_ _231_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__or2_1
XFILLER_12_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_484_ net11 net8 net45 _109_ net13 VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__o41a_1
X_622_ counter\[19\] counter\[18\] _277_ VGND VGND VPWR VPWR _282_ sky130_fd_sc_hd__and3_1
XFILLER_8_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_398_ net22 VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__inv_2
X_467_ _141_ _143_ _144_ _145_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__and4_1
X_536_ counter\[6\] _214_ VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__or2_1
X_605_ counter\[14\] _269_ VGND VGND VPWR VPWR _270_ sky130_fd_sc_hd__nand2_1
Xfanout40 net33 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_0_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_519_ _071_ _099_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__xnor2_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_784_ clknet_2_0__leaf_clk _002_ _045_ VGND VGND VPWR VPWR counter\[11\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_6_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_767_ net43 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__inv_2
XFILLER_21_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_698_ _342_ _343_ _344_ VGND VGND VPWR VPWR _345_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_15_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_552_ _134_ _124_ _147_ _230_ VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__nand4_2
XTAP_TAPCELL_ROW_23_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_483_ counter\[21\] _160_ _161_ _159_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__o211ai_1
XFILLER_12_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_621_ counter\[19\] _279_ VGND VGND VPWR VPWR _281_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_20_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_466_ counter\[25\] _137_ VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__or2_1
X_535_ _099_ _213_ VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__and2_1
X_604_ _269_ net35 _268_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and3b_1
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_397_ counter\[9\] VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout41 net33 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_449_ counter\[29\] _125_ _127_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__a21oi_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_518_ _100_ _196_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_783_ clknet_2_0__leaf_clk _001_ _044_ VGND VGND VPWR VPWR counter\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_6_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_697_ net26 counter\[2\] VGND VGND VPWR VPWR _344_ sky130_fd_sc_hd__xor2_1
X_766_ net43 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_23_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_551_ _139_ _145_ _229_ VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__and3b_1
X_620_ _279_ _280_ net35 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__and3b_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_482_ _154_ _157_ counter\[22\] VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__a21o_1
XFILLER_12_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_3_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_749_ net40 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__inv_2
XFILLER_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_465_ counter\[26\] _142_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__or2_1
X_534_ _069_ _098_ _070_ VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__a21o_1
X_603_ counter\[13\] counter\[12\] counter\[11\] _262_ VGND VGND VPWR VPWR _269_ sky130_fd_sc_hd__and4_1
XFILLER_5_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_396_ counter\[10\] VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__inv_2
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout42 net33 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_4
X_448_ counter\[28\] _117_ _126_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__and3_1
X_517_ net30 net44 net31 VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_0_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_782_ clknet_2_0__leaf_clk _031_ _043_ VGND VGND VPWR VPWR counter\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_696_ counter\[3\] net27 VGND VGND VPWR VPWR _343_ sky130_fd_sc_hd__and2b_1
X_765_ net43 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_550_ counter\[24\] _138_ VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_481_ net14 _153_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_748_ net40 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__inv_2
X_679_ _087_ counter\[17\] counter\[16\] _088_ VGND VGND VPWR VPWR _326_ sky130_fd_sc_hd__o22a_1
X_464_ counter\[26\] _142_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__nand2_1
X_533_ counter\[4\] _209_ _211_ counter\[5\] VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__a22o_1
X_602_ counter\[13\] _267_ VGND VGND VPWR VPWR _268_ sky130_fd_sc_hd__or2_1
X_395_ counter\[12\] VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__inv_2
Xfanout43 net33 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_447_ net39 _111_ _115_ _079_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__a31o_1
X_516_ counter\[9\] _193_ VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_0_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_781_ clknet_2_0__leaf_clk _030_ _042_ VGND VGND VPWR VPWR counter\[8\] sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_10_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_695_ net27 counter\[3\] VGND VGND VPWR VPWR _342_ sky130_fd_sc_hd__and2b_1
X_764_ net43 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_31_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_480_ _113_ _155_ counter\[23\] VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__a21o_1
XFILLER_16_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_747_ net42 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__inv_2
X_678_ _086_ counter\[18\] _324_ VGND VGND VPWR VPWR _325_ sky130_fd_sc_hd__a21bo_1
X_601_ _267_ net35 _266_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and3b_1
X_463_ _080_ _114_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__xnor2_1
X_532_ net28 _098_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_394_ counter\[13\] VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__inv_2
X_446_ _078_ _117_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_0_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_515_ counter\[10\] _192_ _193_ counter\[9\] VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__a22o_1
X_429_ net16 net13 net11 net8 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__or4_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 psc[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_6
XFILLER_19_118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_780_ clknet_2_2__leaf_clk _029_ _041_ VGND VGND VPWR VPWR counter\[7\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_7_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_694_ _070_ counter\[5\] counter\[4\] _069_ VGND VGND VPWR VPWR _341_ sky130_fd_sc_hd__a22o_1
X_763_ net42 VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__inv_2
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_31_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_746_ net42 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__inv_2
X_677_ counter\[19\] net13 VGND VGND VPWR VPWR _324_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_462_ _116_ _140_ counter\[27\] VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__a21o_1
X_531_ counter\[3\] _200_ _209_ counter\[4\] _207_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__o221a_1
X_600_ counter\[12\] counter\[11\] _262_ VGND VGND VPWR VPWR _267_ sky130_fd_sc_hd__and3_1
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_393_ counter\[14\] VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__inv_2
X_729_ _362_ _370_ _375_ _338_ VGND VGND VPWR VPWR _376_ sky130_fd_sc_hd__o31a_1
X_514_ _072_ _100_ VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__xnor2_1
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_445_ _120_ _119_ counter\[31\] _123_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__a31oi_4
XPHY_EDGE_ROW_23_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_428_ net6 net7 _104_ _103_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__or4_4
XFILLER_10_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput2 psc[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_693_ _071_ counter\[6\] VGND VGND VPWR VPWR _340_ sky130_fd_sc_hd__and2_1
X_762_ net41 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__inv_2
XFILLER_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_10_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_745_ net42 VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__inv_2
X_676_ _086_ counter\[18\] VGND VGND VPWR VPWR _323_ sky130_fd_sc_hd__nor2_1
X_461_ net19 _114_ net20 VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__o21ai_1
X_530_ _098_ _208_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__and2b_1
X_392_ net32 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__inv_2
XFILLER_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_659_ _090_ counter\[29\] VGND VGND VPWR VPWR _306_ sky130_fd_sc_hd__and2_1
X_728_ _364_ _374_ _363_ VGND VGND VPWR VPWR _375_ sky130_fd_sc_hd__o21a_1
Xfanout35 _243_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_6
X_444_ _118_ counter\[30\] _122_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__and3_1
X_513_ net2 _101_ VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__xor2_1
XFILLER_24_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_427_ net6 net7 net46 _104_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nor4_4
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 psc[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_761_ net41 VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_17_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_692_ counter\[7\] net31 VGND VGND VPWR VPWR _339_ sky130_fd_sc_hd__nand2b_1
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_744_ net42 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_675_ net13 counter\[19\] VGND VGND VPWR VPWR _322_ sky130_fd_sc_hd__and2b_1
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_460_ counter\[25\] _137_ _138_ counter\[24\] VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__a22o_1
X_391_ net30 VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__inv_2
X_658_ _078_ counter\[28\] VGND VGND VPWR VPWR _305_ sky130_fd_sc_hd__and2_1
XFILLER_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_727_ _359_ _373_ _357_ VGND VGND VPWR VPWR _374_ sky130_fd_sc_hd__a21oi_1
X_589_ _077_ _257_ VGND VGND VPWR VPWR _259_ sky130_fd_sc_hd__nand2_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout36 _243_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_6
XFILLER_1_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_443_ net22 net47 net24 VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__o21ai_1
XFILLER_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_512_ _103_ _190_ VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__and2_1
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 psc[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_426_ _103_ _104_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nor2_1
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_409_ net8 VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__inv_2
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_691_ _333_ _334_ _337_ VGND VGND VPWR VPWR _338_ sky130_fd_sc_hd__nor3_1
XFILLER_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_760_ net41 VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__inv_2
X_743_ net42 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_22_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_674_ _084_ counter\[21\] counter\[20\] _085_ VGND VGND VPWR VPWR _321_ sky130_fd_sc_hd__a22o_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_390_ net29 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__inv_2
X_657_ counter\[31\] _304_ net38 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__o21a_1
X_588_ net35 _257_ _258_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__and3_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_726_ _371_ _372_ VGND VGND VPWR VPWR _373_ sky130_fd_sc_hd__nand2_1
Xfanout37 _243_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_6
XFILLER_13_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_442_ _119_ _120_ counter\[31\] VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_511_ net2 _101_ net3 VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_709_ net6 _074_ _075_ net5 VGND VGND VPWR VPWR _356_ sky130_fd_sc_hd__o22a_1
XFILLER_24_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 psc[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_425_ net5 net4 VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_27_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_408_ net9 VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_690_ _317_ _320_ _335_ _336_ VGND VGND VPWR VPWR _337_ sky130_fd_sc_hd__or4b_1
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput30 psc[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_22_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_742_ net42 VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__inv_2
X_673_ _083_ counter\[22\] VGND VGND VPWR VPWR _320_ sky130_fd_sc_hd__and2_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_656_ _304_ net38 _303_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__and3b_1
Xclone11 _243_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
X_587_ counter\[8\] _255_ VGND VGND VPWR VPWR _258_ sky130_fd_sc_hd__or2_1
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_725_ net3 _076_ _355_ _360_ _358_ VGND VGND VPWR VPWR _372_ sky130_fd_sc_hd__a221o_1
Xfanout38 _243_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_6
X_441_ net22 net24 net25 net48 VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__or4_4
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_510_ counter\[13\] _185_ _188_ counter\[12\] VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__a22o_1
X_639_ counter\[24\] _290_ counter\[25\] VGND VGND VPWR VPWR _293_ sky130_fd_sc_hd__a21o_1
X_708_ net65 _072_ net2 _077_ VGND VGND VPWR VPWR _355_ sky130_fd_sc_hd__a2bb2o_4
XTAP_TAPCELL_ROW_1_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_424_ net30 net3 _102_ _099_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__or4_4
XFILLER_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput6 psc[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_407_ net10 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_25_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput20 psc[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 psc[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_22_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_741_ net42 VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__inv_2
X_672_ _083_ counter\[22\] VGND VGND VPWR VPWR _319_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_31_Left_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_724_ _358_ _361_ VGND VGND VPWR VPWR _371_ sky130_fd_sc_hd__nand2b_1
X_655_ _092_ _302_ VGND VGND VPWR VPWR _304_ sky130_fd_sc_hd__nor2_1
X_586_ net63 _255_ VGND VGND VPWR VPWR _257_ sky130_fd_sc_hd__nand2_1
X_440_ net22 net24 _117_ net25 VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o31ai_4
X_569_ counter\[0\] counter\[1\] counter\[2\] VGND VGND VPWR VPWR _246_ sky130_fd_sc_hd__a21o_1
X_638_ net54 _291_ _292_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__and3_1
X_707_ _340_ _353_ _339_ VGND VGND VPWR VPWR _354_ sky130_fd_sc_hd__o21ai_1
X_423_ net2 net32 net31 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__or3_1
Xinput7 psc[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_28_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_406_ net11 VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__inv_2
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput21 psc[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput32 psc[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xinput10 psc[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
X_740_ net42 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__inv_2
X_671_ _082_ counter\[23\] VGND VGND VPWR VPWR _318_ sky130_fd_sc_hd__nor2_1
XFILLER_4_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_654_ _092_ _302_ VGND VGND VPWR VPWR _303_ sky130_fd_sc_hd__nand2_1
X_723_ _368_ _369_ _354_ VGND VGND VPWR VPWR _370_ sky130_fd_sc_hd__and3b_1
X_585_ _255_ _256_ net35 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__and3b_1
XFILLER_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_637_ counter\[24\] _290_ VGND VGND VPWR VPWR _292_ sky130_fd_sc_hd__or2_1
X_706_ _071_ counter\[6\] counter\[5\] _070_ _352_ VGND VGND VPWR VPWR _353_ sky130_fd_sc_hd__o221a_1
X_568_ counter\[0\] counter\[1\] counter\[2\] VGND VGND VPWR VPWR _245_ sky130_fd_sc_hd__and3_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_499_ _175_ _177_ _172_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__and3b_1
X_422_ net30 net32 net31 _099_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__or4_1
Xinput8 psc[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_405_ net14 VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__inv_2
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput22 psc[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_1
Xinput33 rst VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 psc[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_670_ _082_ counter\[23\] VGND VGND VPWR VPWR _317_ sky130_fd_sc_hd__and2_1
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_799_ clknet_2_3__leaf_clk _018_ _060_ VGND VGND VPWR VPWR counter\[26\] sky130_fd_sc_hd__dfrtp_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_653_ net38 _301_ _302_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__and3_1
X_722_ net31 counter\[7\] VGND VGND VPWR VPWR _369_ sky130_fd_sc_hd__nand2b_1
X_584_ counter\[7\] _253_ VGND VGND VPWR VPWR _256_ sky130_fd_sc_hd__or2_1
XFILLER_4_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_567_ net37 _204_ _244_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__and3_1
X_705_ _348_ _349_ _351_ _341_ VGND VGND VPWR VPWR _352_ sky130_fd_sc_hd__a31o_1
X_636_ counter\[24\] _290_ VGND VGND VPWR VPWR _291_ sky130_fd_sc_hd__nand2_1
X_498_ counter\[17\] _174_ _176_ counter\[16\] VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__a22o_1
X_421_ net30 net31 _099_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__or3_1
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_619_ counter\[18\] _277_ VGND VGND VPWR VPWR _280_ sky130_fd_sc_hd__or2_1
Xinput9 psc[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_1
X_404_ net15 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__inv_2
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_6_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput23 psc[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 psc[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_6
XFILLER_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_798_ clknet_2_3__leaf_clk _017_ _059_ VGND VGND VPWR VPWR counter\[25\] sky130_fd_sc_hd__dfrtp_1
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_652_ counter\[29\] _299_ VGND VGND VPWR VPWR _302_ sky130_fd_sc_hd__nand2_1
X_583_ counter\[7\] _253_ VGND VGND VPWR VPWR _255_ sky130_fd_sc_hd__and2_1
X_721_ _361_ _362_ _367_ _365_ VGND VGND VPWR VPWR _368_ sky130_fd_sc_hd__or4_4
XPHY_EDGE_ROW_9_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_566_ counter\[0\] counter\[1\] VGND VGND VPWR VPWR _244_ sky130_fd_sc_hd__or2_1
X_704_ _343_ _350_ VGND VGND VPWR VPWR _351_ sky130_fd_sc_hd__nor2_1
X_635_ _290_ net54 _289_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__and3b_1
XFILLER_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_497_ net8 _106_ VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__xnor2_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_420_ net28 net27 _097_ net29 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__or4_4
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_549_ _158_ _159_ VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__nand2_1
X_618_ counter\[18\] _277_ VGND VGND VPWR VPWR _279_ sky130_fd_sc_hd__and2_1
X_403_ net16 VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__inv_2
XFILLER_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_22_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap39 _106_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
Xinput24 psc[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 psc[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_21_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_797_ clknet_2_3__leaf_clk _016_ _058_ VGND VGND VPWR VPWR counter\[24\] sky130_fd_sc_hd__dfrtp_2
X_651_ counter\[29\] _299_ VGND VGND VPWR VPWR _301_ sky130_fd_sc_hd__or2_1
X_582_ _253_ _254_ net37 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and3b_1
X_720_ _355_ _357_ _364_ _366_ VGND VGND VPWR VPWR _367_ sky130_fd_sc_hd__or4_4
X_565_ _066_ net54 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and2_1
XFILLER_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_703_ _069_ counter\[4\] VGND VGND VPWR VPWR _350_ sky130_fd_sc_hd__nor2_1
X_634_ counter\[23\] counter\[22\] counter\[21\] _283_ VGND VGND VPWR VPWR _290_ sky130_fd_sc_hd__and4_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_496_ counter\[17\] _174_ VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__nor2_1
XFILLER_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_479_ counter\[22\] _154_ _157_ _156_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__a31o_1
X_548_ _158_ _162_ _165_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__or3_1
X_617_ counter\[17\] _274_ _278_ net35 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__o211a_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_402_ net17 VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__inv_2
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput25 psc[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_1
Xinput14 psc[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_796_ clknet_2_3__leaf_clk _015_ _057_ VGND VGND VPWR VPWR counter\[23\] sky130_fd_sc_hd__dfrtp_1
X_650_ _299_ _300_ net38 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__and3b_1
X_581_ counter\[6\] _251_ VGND VGND VPWR VPWR _254_ sky130_fd_sc_hd__or2_1
X_779_ clknet_2_2__leaf_clk _028_ _040_ VGND VGND VPWR VPWR counter\[6\] sky130_fd_sc_hd__dfrtp_1
X_702_ counter\[2\] _342_ net26 VGND VGND VPWR VPWR _349_ sky130_fd_sc_hd__or3b_1
X_564_ _232_ _242_ _151_ _241_ VGND VGND VPWR VPWR _243_ sky130_fd_sc_hd__o211a_4
X_633_ counter\[23\] _287_ VGND VGND VPWR VPWR _289_ sky130_fd_sc_hd__or2_1
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_495_ _168_ _173_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__and2_4
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_478_ _085_ _153_ _084_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__a21o_1
X_547_ _158_ _162_ _166_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__or3_1
X_616_ _277_ VGND VGND VPWR VPWR _278_ sky130_fd_sc_hd__inv_2
X_401_ net18 VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__inv_2
XFILLER_2_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput26 psc[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
Xinput15 psc[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_21_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_146 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_795_ clknet_2_1__leaf_clk _014_ _056_ VGND VGND VPWR VPWR counter\[22\] sky130_fd_sc_hd__dfrtp_1
X_580_ counter\[6\] counter\[5\] counter\[4\] _247_ VGND VGND VPWR VPWR _253_ sky130_fd_sc_hd__and4_1
X_778_ clknet_2_2__leaf_clk _027_ _039_ VGND VGND VPWR VPWR counter\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_28_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_701_ _346_ _347_ _345_ VGND VGND VPWR VPWR _348_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_632_ _287_ _288_ net36 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__and3b_1
X_563_ _179_ _226_ _227_ _228_ VGND VGND VPWR VPWR _242_ sky130_fd_sc_hd__o211a_1
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_494_ _089_ net39 _088_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__a21o_1
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_477_ counter\[23\] _113_ _155_ VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__and3_1
X_615_ counter\[15\] counter\[14\] _269_ _276_ VGND VGND VPWR VPWR _277_ sky130_fd_sc_hd__and4_1
X_546_ counter\[16\] _176_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__nor2_1
XFILLER_25_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_400_ net19 VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__inv_2
XFILLER_18_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_529_ net27 _097_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_19_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_26_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput27 psc[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_16_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput16 psc[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_1
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_794_ clknet_2_1__leaf_clk _013_ _055_ VGND VGND VPWR VPWR counter\[21\] sky130_fd_sc_hd__dfrtp_4
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_29_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_777_ clknet_2_2__leaf_clk _026_ _038_ VGND VGND VPWR VPWR counter\[4\] sky130_fd_sc_hd__dfrtp_4
XPHY_EDGE_ROW_13_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_700_ _066_ net12 counter\[1\] _068_ VGND VGND VPWR VPWR _347_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_562_ _148_ _231_ _237_ _240_ VGND VGND VPWR VPWR _241_ sky130_fd_sc_hd__or4_4
X_631_ counter\[21\] _283_ counter\[22\] VGND VGND VPWR VPWR _288_ sky130_fd_sc_hd__a21o_1
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_493_ counter\[19\] _167_ _169_ counter\[18\] VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__o22a_1
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_476_ _084_ _085_ _153_ _083_ VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__a31o_1
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_614_ counter\[17\] counter\[16\] VGND VGND VPWR VPWR _276_ sky130_fd_sc_hd__and2_1
X_545_ _218_ _222_ _223_ _220_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__a31o_1
XFILLER_25_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_528_ counter\[3\] _200_ _202_ _206_ _203_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_19_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_459_ _082_ _113_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__xnor2_1
XFILLER_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 psc[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
Xinput28 psc[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_793_ clknet_2_1__leaf_clk _012_ _054_ VGND VGND VPWR VPWR counter\[20\] sky130_fd_sc_hd__dfrtp_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_776_ clknet_2_3__leaf_clk _025_ _037_ VGND VGND VPWR VPWR counter\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_30_Left_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_630_ counter\[22\] counter\[21\] _283_ VGND VGND VPWR VPWR _287_ sky130_fd_sc_hd__and3_1
X_561_ _158_ _162_ _166_ _239_ VGND VGND VPWR VPWR _240_ sky130_fd_sc_hd__or4_4
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_492_ counter\[19\] _167_ _170_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__o21a_1
X_759_ net41 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__inv_2
X_613_ _274_ _275_ net36 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__and3b_1
X_544_ _216_ _217_ _194_ VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__o21ba_1
X_475_ net15 net14 _153_ VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__or3b_1
XFILLER_26_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_527_ _095_ _205_ _204_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__a21bo_1
X_458_ _114_ _136_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__and2_1
X_389_ net28 VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__inv_2
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 psc[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_1
Xinput29 psc[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_792_ clknet_2_1__leaf_clk _010_ _053_ VGND VGND VPWR VPWR counter\[19\] sky130_fd_sc_hd__dfrtp_2
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_775_ clknet_2_2__leaf_clk _022_ _036_ VGND VGND VPWR VPWR counter\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_560_ _175_ _177_ _238_ _172_ VGND VGND VPWR VPWR _239_ sky130_fd_sc_hd__or4b_4
X_491_ counter\[19\] _167_ _169_ counter\[18\] VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_689_ _084_ counter\[21\] counter\[20\] _085_ VGND VGND VPWR VPWR _336_ sky130_fd_sc_hd__o22a_1
X_758_ net41 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__inv_2
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_543_ net62 _197_ _198_ counter\[7\] _221_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__o221a_1
X_474_ _109_ _089_ _106_ _112_ VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__and4b_1
X_612_ counter\[16\] _273_ VGND VGND VPWR VPWR _275_ sky130_fd_sc_hd__or2_1
XFILLER_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_27_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_526_ net1 _066_ net12 _067_ VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__o211ai_1
XFILLER_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_388_ net23 VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__inv_2
XFILLER_23_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_457_ _082_ net39 _111_ _081_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__a31o_1
Xinput19 psc[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_1
XFILLER_14_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_509_ _184_ _187_ VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__and2_1
X_791_ clknet_2_1__leaf_clk _009_ _052_ VGND VGND VPWR VPWR counter\[18\] sky130_fd_sc_hd__dfrtp_4
XFILLER_6_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_774_ clknet_2_2__leaf_clk _011_ _035_ VGND VGND VPWR VPWR counter\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_490_ net10 _168_ _152_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_17_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_757_ net40 VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__inv_2
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_688_ _088_ counter\[16\] _322_ _323_ _327_ VGND VGND VPWR VPWR _335_ sky130_fd_sc_hd__a2111o_1
X_542_ net62 _197_ _193_ counter\[9\] VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__o2bb2a_1
X_611_ counter\[16\] _273_ VGND VGND VPWR VPWR _274_ sky130_fd_sc_hd__and2_1
X_473_ _109_ _089_ _106_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__and3b_1
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer20 net62 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_525_ counter\[0\] counter\[1\] VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__nand2_1
X_387_ counter\[1\] VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__inv_2
X_456_ _124_ _134_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__and2_1
XFILLER_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_439_ net22 net24 _117_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__or3_4
X_508_ net4 _103_ VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_30_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_790_ clknet_2_1__leaf_clk _008_ _051_ VGND VGND VPWR VPWR counter\[17\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_5_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_773_ clknet_2_2__leaf_clk _000_ _034_ VGND VGND VPWR VPWR counter\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_687_ _325_ _326_ VGND VGND VPWR VPWR _334_ sky130_fd_sc_hd__nand2b_1
X_756_ net40 VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_8_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_472_ _135_ _150_ _121_ _131_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__o2bb2a_1
X_610_ _273_ net36 _272_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and3b_1
X_541_ counter\[11\] _191_ _218_ _219_ VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__a22o_1
X_739_ _368_ _384_ _385_ _380_ _377_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__o32a_1
XFILLER_26_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer21 net62 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd1_1
X_386_ counter\[0\] VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__inv_2
X_455_ _121_ _129_ _133_ _130_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__nor4_4
X_524_ counter\[2\] _096_ _201_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__and3_1
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_438_ net21 _110_ net45 _115_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__or4b_4
Xrebuffer1 _099_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_11_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_507_ counter\[14\] _182_ _185_ counter\[13\] VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__o22a_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_772_ clknet_2_2__leaf_clk _032_ _033_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_755_ net40 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__inv_2
X_686_ _318_ _321_ _319_ VGND VGND VPWR VPWR _333_ sky130_fd_sc_hd__or3b_1
XTAP_TAPCELL_ROW_5_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_471_ _139_ _146_ _148_ _149_ VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__a211o_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_540_ net64 _195_ _197_ _194_ VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__a31o_1
X_669_ _310_ _312_ _313_ _315_ VGND VGND VPWR VPWR _316_ sky130_fd_sc_hd__and4_1
X_738_ _316_ _338_ VGND VGND VPWR VPWR _385_ sky130_fd_sc_hd__nand2_1
Xrebuffer22 counter\[8\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_6
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_454_ counter\[29\] _125_ _127_ _132_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__a211o_1
X_523_ _096_ _201_ counter\[2\] VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__a21o_1
XFILLER_17_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ net20 net19 _114_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_15_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_506_ net5 _184_ _105_ VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer2 _107_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_771_ net43 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__inv_2
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_685_ _317_ _331_ VGND VGND VPWR VPWR _332_ sky130_fd_sc_hd__nor2_1
X_754_ net40 VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_737_ _382_ _383_ _346_ VGND VGND VPWR VPWR _384_ sky130_fd_sc_hd__or3b_1
X_470_ counter\[26\] _141_ _142_ VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__and3_1
X_668_ _314_ VGND VGND VPWR VPWR _315_ sky130_fd_sc_hd__inv_2
X_599_ counter\[12\] _265_ VGND VGND VPWR VPWR _266_ sky130_fd_sc_hd__or2_1
XFILLER_26_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_522_ net23 _095_ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__nand2_1
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_453_ _117_ _126_ counter\[28\] VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__a21oi_1
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_436_ net20 _080_ _081_ _082_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__and4b_1
XTAP_TAPCELL_ROW_15_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_505_ net4 _103_ VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__or2_1
Xrebuffer3 _103_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
XFILLER_9_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_419_ net27 _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__nor2_1
X_770_ net43 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__inv_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_684_ _082_ counter\[23\] _320_ _330_ _319_ VGND VGND VPWR VPWR _331_ sky130_fd_sc_hd__o221a_1
X_753_ net40 VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__inv_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_736_ _066_ net12 _340_ _345_ _350_ VGND VGND VPWR VPWR _383_ sky130_fd_sc_hd__a2111o_1
XFILLER_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_667_ net20 _094_ counter\[25\] _080_ VGND VGND VPWR VPWR _314_ sky130_fd_sc_hd__a2bb2o_1
X_598_ _265_ net35 _264_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__and3b_1
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_452_ _128_ _129_ _130_ _124_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__o31a_1
X_521_ _097_ _199_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__and2_1
XFILLER_31_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_719_ _360_ _363_ VGND VGND VPWR VPWR _366_ sky130_fd_sc_hd__nand2_1
XFILLER_22_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer4 net48 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_435_ net18 net17 net45 _110_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__or4_4
XTAP_TAPCELL_ROW_15_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_504_ counter\[15\] _181_ _182_ counter\[14\] VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__a22o_1
XFILLER_22_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_418_ net1 net12 net26 net23 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__or4_4
XPHY_EDGE_ROW_25_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_683_ _084_ counter\[21\] _321_ _329_ VGND VGND VPWR VPWR _330_ sky130_fd_sc_hd__o22a_1
X_752_ net40 VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__inv_2
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_804_ clknet_2_3__leaf_clk _024_ _065_ VGND VGND VPWR VPWR counter\[31\] sky130_fd_sc_hd__dfrtp_1
XFILLER_29_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_735_ _341_ _347_ _381_ _339_ VGND VGND VPWR VPWR _382_ sky130_fd_sc_hd__or4bb_1
X_666_ _080_ counter\[25\] counter\[24\] _081_ VGND VGND VPWR VPWR _313_ sky130_fd_sc_hd__o22a_1
X_597_ counter\[11\] _262_ VGND VGND VPWR VPWR _265_ sky130_fd_sc_hd__and2_1
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_520_ net26 _096_ VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__nand2_1
X_451_ _118_ _122_ counter\[30\] VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__a21oi_1
X_649_ counter\[27\] _295_ counter\[28\] VGND VGND VPWR VPWR _300_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_18_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_718_ net3 _076_ net65 _072_ _358_ VGND VGND VPWR VPWR _365_ sky130_fd_sc_hd__a221o_1
XFILLER_16_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_434_ net39 _111_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__nand2_1
X_503_ net6 _105_ VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__xnor2_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xrebuffer5 _117_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_0_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_417_ net1 net12 net23 VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__or3_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_682_ _085_ counter\[20\] _322_ _328_ _324_ VGND VGND VPWR VPWR _329_ sky130_fd_sc_hd__o221a_1
X_751_ net40 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_803_ clknet_2_3__leaf_clk _023_ _064_ VGND VGND VPWR VPWR counter\[30\] sky130_fd_sc_hd__dfrtp_2
XFILLER_29_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_665_ _081_ counter\[24\] _311_ VGND VGND VPWR VPWR _312_ sky130_fd_sc_hd__a21oi_1
X_734_ _071_ counter\[6\] counter\[5\] _070_ _369_ VGND VGND VPWR VPWR _381_ sky130_fd_sc_hd__o221a_1
X_596_ counter\[11\] _262_ VGND VGND VPWR VPWR _264_ sky130_fd_sc_hd__or2_1
XFILLER_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_450_ counter\[29\] _125_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__nor2_1
X_648_ counter\[28\] counter\[27\] _295_ VGND VGND VPWR VPWR _299_ sky130_fd_sc_hd__and3_1
X_579_ _251_ _252_ net37 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and3b_1
XFILLER_16_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_717_ net7 _073_ _074_ net6 VGND VGND VPWR VPWR _364_ sky130_fd_sc_hd__a22o_1
XFILLER_26_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_433_ net13 net11 VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__nor2_1
X_502_ _106_ _180_ VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__nor2_1
XFILLER_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_416_ net1 net12 VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__or2_1
XFILLER_12_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_750_ net40 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__inv_2
X_681_ _325_ _326_ _327_ counter\[18\] _086_ VGND VGND VPWR VPWR _328_ sky130_fd_sc_hd__o32a_1
XFILLER_22_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_802_ clknet_2_3__leaf_clk _021_ _063_ VGND VGND VPWR VPWR counter\[29\] sky130_fd_sc_hd__dfrtp_2
X_733_ _310_ _378_ _379_ _307_ VGND VGND VPWR VPWR _380_ sky130_fd_sc_hd__a22o_1
X_664_ net21 _093_ _094_ net20 VGND VGND VPWR VPWR _311_ sky130_fd_sc_hd__a22o_1
X_595_ _262_ _263_ net35 VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__and3b_1
XFILLER_6_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_647_ net54 _297_ _298_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__and3_1
X_578_ counter\[4\] _247_ counter\[5\] VGND VGND VPWR VPWR _252_ sky130_fd_sc_hd__a21o_1
XFILLER_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_716_ counter\[15\] _089_ _073_ net7 VGND VGND VPWR VPWR _363_ sky130_fd_sc_hd__o2bb2a_1
.ends

