magic
tech sky130A
magscale 1 2
timestamp 1729848072
<< error_p >>
rect -29 525 29 531
rect -29 491 -17 525
rect -29 485 29 491
<< nwell >>
rect -112 -578 112 544
<< pmos >>
rect -18 -516 18 444
<< pdiff >>
rect -76 432 -18 444
rect -76 -504 -64 432
rect -30 -504 -18 432
rect -76 -516 -18 -504
rect 18 432 76 444
rect 18 -504 30 432
rect 64 -504 76 432
rect 18 -516 76 -504
<< pdiffc >>
rect -64 -504 -30 432
rect 30 -504 64 432
<< poly >>
rect -33 525 33 541
rect -33 491 -17 525
rect 17 491 33 525
rect -33 475 33 491
rect -18 444 18 475
rect -18 -542 18 -516
<< polycont >>
rect -17 491 17 525
<< locali >>
rect -33 491 -17 525
rect 17 491 33 525
rect -64 432 -30 448
rect -64 -520 -30 -504
rect 30 432 64 448
rect 30 -520 64 -504
<< viali >>
rect -17 491 17 525
rect -64 -504 -30 432
rect 30 -504 64 432
<< metal1 >>
rect -29 525 29 531
rect -29 491 -17 525
rect 17 491 29 525
rect -29 485 29 491
rect -70 432 -24 444
rect -70 -504 -64 432
rect -30 -504 -24 432
rect -70 -516 -24 -504
rect 24 432 70 444
rect 24 -504 30 432
rect 64 -504 70 432
rect 24 -516 70 -504
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.8 l 0.18 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
