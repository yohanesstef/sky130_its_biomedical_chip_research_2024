VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO freq_psc
  CLASS BLOCK ;
  FOREIGN freq_psc ;
  ORIGIN 0.000 0.000 ;
  SIZE 83.030 BY 93.750 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 81.840 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 81.840 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END clk
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END out
  PIN psc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 27.240 83.030 27.840 ;
    END
  END psc[0]
  PIN psc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 89.750 55.110 93.750 ;
    END
  END psc[10]
  PIN psc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 89.750 58.330 93.750 ;
    END
  END psc[11]
  PIN psc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 89.750 42.230 93.750 ;
    END
  END psc[12]
  PIN psc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 89.750 45.450 93.750 ;
    END
  END psc[13]
  PIN psc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 89.750 51.890 93.750 ;
    END
  END psc[14]
  PIN psc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 89.750 48.670 93.750 ;
    END
  END psc[15]
  PIN psc[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 51.040 83.030 51.640 ;
    END
  END psc[16]
  PIN psc[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 44.240 83.030 44.840 ;
    END
  END psc[17]
  PIN psc[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END psc[18]
  PIN psc[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END psc[19]
  PIN psc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 34.040 83.030 34.640 ;
    END
  END psc[1]
  PIN psc[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END psc[20]
  PIN psc[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END psc[21]
  PIN psc[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END psc[22]
  PIN psc[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END psc[23]
  PIN psc[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END psc[24]
  PIN psc[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END psc[25]
  PIN psc[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END psc[26]
  PIN psc[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END psc[27]
  PIN psc[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END psc[28]
  PIN psc[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END psc[29]
  PIN psc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 30.640 83.030 31.240 ;
    END
  END psc[2]
  PIN psc[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END psc[30]
  PIN psc[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END psc[31]
  PIN psc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 37.440 83.030 38.040 ;
    END
  END psc[3]
  PIN psc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 40.840 83.030 41.440 ;
    END
  END psc[4]
  PIN psc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 47.640 83.030 48.240 ;
    END
  END psc[5]
  PIN psc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 54.440 83.030 55.040 ;
    END
  END psc[6]
  PIN psc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 57.840 83.030 58.440 ;
    END
  END psc[7]
  PIN psc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 61.240 83.030 61.840 ;
    END
  END psc[8]
  PIN psc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 64.640 83.030 65.240 ;
    END
  END psc[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 79.030 17.040 83.030 17.640 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 77.470 81.685 ;
      LAYER li1 ;
        RECT 5.520 10.795 77.280 81.685 ;
      LAYER met1 ;
        RECT 4.210 10.640 77.280 81.840 ;
      LAYER met2 ;
        RECT 4.230 89.470 41.670 89.750 ;
        RECT 42.510 89.470 44.890 89.750 ;
        RECT 45.730 89.470 48.110 89.750 ;
        RECT 48.950 89.470 51.330 89.750 ;
        RECT 52.170 89.470 54.550 89.750 ;
        RECT 55.390 89.470 57.770 89.750 ;
        RECT 58.610 89.470 76.270 89.750 ;
        RECT 4.230 4.280 76.270 89.470 ;
        RECT 4.230 4.000 19.130 4.280 ;
        RECT 19.970 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 76.270 4.280 ;
      LAYER met3 ;
        RECT 3.990 75.840 79.030 81.765 ;
        RECT 4.400 74.440 79.030 75.840 ;
        RECT 3.990 65.640 79.030 74.440 ;
        RECT 4.400 64.240 78.630 65.640 ;
        RECT 3.990 62.240 79.030 64.240 ;
        RECT 4.400 60.840 78.630 62.240 ;
        RECT 3.990 58.840 79.030 60.840 ;
        RECT 4.400 57.440 78.630 58.840 ;
        RECT 3.990 55.440 79.030 57.440 ;
        RECT 4.400 54.040 78.630 55.440 ;
        RECT 3.990 52.040 79.030 54.040 ;
        RECT 4.400 50.640 78.630 52.040 ;
        RECT 3.990 48.640 79.030 50.640 ;
        RECT 4.400 47.240 78.630 48.640 ;
        RECT 3.990 45.240 79.030 47.240 ;
        RECT 4.400 43.840 78.630 45.240 ;
        RECT 3.990 41.840 79.030 43.840 ;
        RECT 4.400 40.440 78.630 41.840 ;
        RECT 3.990 38.440 79.030 40.440 ;
        RECT 4.400 37.040 78.630 38.440 ;
        RECT 3.990 35.040 79.030 37.040 ;
        RECT 3.990 33.640 78.630 35.040 ;
        RECT 3.990 31.640 79.030 33.640 ;
        RECT 4.400 30.240 78.630 31.640 ;
        RECT 3.990 28.240 79.030 30.240 ;
        RECT 3.990 26.840 78.630 28.240 ;
        RECT 3.990 18.040 79.030 26.840 ;
        RECT 3.990 16.640 78.630 18.040 ;
        RECT 3.990 10.715 79.030 16.640 ;
  END
END freq_psc
END LIBRARY

