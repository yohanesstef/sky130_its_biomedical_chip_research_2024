magic
tech sky130A
magscale 1 2
timestamp 1730525416
<< nwell >>
rect -214 -350 214 350
<< pmos >>
rect -120 -250 120 250
<< pdiff >>
rect -178 238 -120 250
rect -178 -238 -166 238
rect -132 -238 -120 238
rect -178 -250 -120 -238
rect 120 238 178 250
rect 120 -238 132 238
rect 166 -238 178 238
rect 120 -250 178 -238
<< pdiffc >>
rect -166 -238 -132 238
rect 132 -238 166 238
<< poly >>
rect -120 331 120 347
rect -120 297 -104 331
rect 104 297 120 331
rect -120 250 120 297
rect -120 -297 120 -250
rect -120 -331 -104 -297
rect 104 -331 120 -297
rect -120 -347 120 -331
<< polycont >>
rect -104 297 104 331
rect -104 -331 104 -297
<< locali >>
rect -120 297 -104 331
rect 104 297 120 331
rect -166 238 -132 254
rect -166 -254 -132 -238
rect 132 238 166 254
rect 132 -254 166 -238
rect -120 -331 -104 -297
rect 104 -331 120 -297
<< viali >>
rect -52 297 52 331
rect -166 -238 -132 238
rect 132 -238 166 238
rect -52 -331 52 -297
<< metal1 >>
rect -64 331 64 337
rect -64 297 -52 331
rect 52 297 64 331
rect -64 291 64 297
rect -172 238 -126 250
rect -172 -238 -166 238
rect -132 -238 -126 238
rect -172 -250 -126 -238
rect 126 238 172 250
rect 126 -238 132 238
rect 166 -238 172 238
rect 126 -250 172 -238
rect -64 -297 64 -291
rect -64 -331 -52 -297
rect 52 -331 64 -297
rect -64 -337 64 -331
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 50 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
