magic
tech sky130A
magscale 1 2
timestamp 1730521008
<< nwell >>
rect -109 -348 109 314
<< pmos >>
rect -15 -286 15 214
<< pdiff >>
rect -73 202 -15 214
rect -73 -274 -61 202
rect -27 -274 -15 202
rect -73 -286 -15 -274
rect 15 202 73 214
rect 15 -274 27 202
rect 61 -274 73 202
rect 15 -286 73 -274
<< pdiffc >>
rect -61 -274 -27 202
rect 27 -274 61 202
<< poly >>
rect -33 295 33 311
rect -33 261 -17 295
rect 17 261 33 295
rect -33 245 33 261
rect -15 214 15 245
rect -15 -312 15 -286
<< polycont >>
rect -17 261 17 295
<< locali >>
rect -33 261 -17 295
rect 17 261 33 295
rect -61 202 -27 218
rect -61 -290 -27 -274
rect 27 202 61 218
rect 27 -290 61 -274
<< viali >>
rect -61 -274 -27 202
rect 27 -274 61 202
<< metal1 >>
rect -67 202 -21 214
rect -67 -274 -61 202
rect -27 -274 -21 202
rect -67 -286 -21 -274
rect 21 202 67 214
rect 21 -274 27 202
rect 61 -274 67 202
rect 21 -286 67 -274
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
