* NGSPICE file created from clk_int_div.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtp_1 abstract view
.subckt sky130_fd_sc_hd__dlxtp_1 D GATE VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd1_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd1_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s4s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s4s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt clk_int_div VGND VPWR clk_i clk_o cycl_count_o[0] cycl_count_o[1] cycl_count_o[2]
+ cycl_count_o[3] cycl_count_o[4] cycl_count_o[5] cycl_count_o[6] cycl_count_o[7]
+ div_i[0] div_i[1] div_i[2] div_i[3] div_i[4] div_i[5] div_i[6] div_i[7] div_ready_o
+ div_valid_i en_i rst_ni test_mode_en_i
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_294_ net35 _013_ net32 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_2
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_277_ net5 div_q\[3\] net24 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__mux2_1
X_200_ even_clk _051_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__xnor2_1
XFILLER_2_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput20 net20 VGND VGND VPWR VPWR cycl_count_o[5] sky130_fd_sc_hd__buf_2
XFILLER_3_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_293_ net35 _012_ net32 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_2
X_276_ net4 div_q\[2\] net24 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__mux2_1
XFILLER_5_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ net15 net16 net17 net18 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__a31o_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput21 net21 VGND VGND VPWR VPWR cycl_count_o[6] sky130_fd_sc_hd__buf_2
XFILLER_22_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_292_ net35 _011_ net32 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_4
XFILLER_3_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_275_ net3 net27 net24 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__mux2_1
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_258_ _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__inv_2
X_189_ div_q\[7\] net9 VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__or2_4
XTAP_TAPCELL_ROW_5_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput22 net22 VGND VGND VPWR VPWR cycl_count_o[7] sky130_fd_sc_hd__buf_2
XFILLER_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_291_ net33 _010_ net30 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_4
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_19_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_274_ div_q\[0\] net24 _108_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_4_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_257_ net15 net16 net17 net18 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__and4_1
XFILLER_9_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_188_ net6 net26 VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_5_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput23 net23 VGND VGND VPWR VPWR div_ready_o sky130_fd_sc_hd__buf_6
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ net34 _009_ net31 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_4
X_273_ _131_ _033_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nor2_1
XFILLER_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_20_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_256_ _093_ _095_ _096_ _091_ net17 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__a32o_1
X_187_ net3 net27 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__xor2_1
X_308_ _000_ _001_ VGND VGND VPWR VPWR i_clk_gate.clk_en sky130_fd_sc_hd__dlxtp_1
XFILLER_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_239_ div_q\[1\] net29 VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__or2_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_272_ net22 _091_ _093_ _107_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a22o_1
XFILLER_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_255_ net29 net16 net17 VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__nand3_1
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ _035_ _036_ _038_ _037_ _034_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__a221o_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_307_ net34 _025_ net31 VGND VGND VPWR VPWR i_clk_mux.clk_sel_i sky130_fd_sc_hd__dfrtp_1
X_169_ net28 net27 VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__xor2_1
X_238_ net27 net29 VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nand2_1
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput14 net14 VGND VGND VPWR VPWR clk_o sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_21_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_271_ net22 _105_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__xnor2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_254_ net29 net16 net17 VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__a21o_1
X_185_ net38 div_q\[6\] VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nand2_1
X_306_ net34 gate_en_d net31 VGND VGND VPWR VPWR gate_en_q sky130_fd_sc_hd__dfrtp_1
X_237_ _122_ _128_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__nand2_1
X_168_ _135_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__inv_2
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_6_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput15 net29 VGND VGND VPWR VPWR cycl_count_o[0] sky130_fd_sc_hd__buf_2
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_16_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_270_ _093_ _105_ _106_ _091_ net21 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__a32o_1
X_253_ _087_ _093_ _094_ _091_ net16 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__a32o_1
X_184_ div_q\[6\] net8 VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__or2_4
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_305_ net34 _024_ net31 VGND VGND VPWR VPWR clk_div_bypass_en_q sky130_fd_sc_hd__dfstp_1
X_236_ net24 _080_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nand2_1
X_167_ clk_div_bypass_en_q net24 _133_ _134_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__and4b_1
X_219_ net28 net29 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_11_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR cycl_count_o[1] sky130_fd_sc_hd__buf_2
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_252_ net15 net16 VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__nand2_1
X_183_ net4 div_q\[2\] VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2_1
X_304_ net34 _023_ net31 VGND VGND VPWR VPWR div_q\[7\] sky130_fd_sc_hd__dfrtp_4
X_235_ _078_ _079_ _134_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__a21o_1
XFILLER_20_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_166_ clk_gate_state_q\[0\] clk_gate_state_q\[1\] VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__nand2b_1
X_218_ div_q\[3\] net18 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__xor2_1
X_149_ net25 _110_ _111_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__o21ba_1
Xoutput17 net17 VGND VGND VPWR VPWR cycl_count_o[2] sky130_fd_sc_hd__buf_2
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_251_ _093_ _091_ net29 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__mux2_1
Xfanout30 net31 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_4
X_182_ net4 div_q\[2\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__or2_4
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_165_ gate_is_open_q clk_gate_state_q\[0\] net10 net11 VGND VGND VPWR VPWR _133_
+ sky130_fd_sc_hd__or4_1
XFILLER_1_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_303_ net33 _022_ net30 VGND VGND VPWR VPWR div_q\[6\] sky130_fd_sc_hd__dfrtp_2
X_234_ _061_ _072_ _073_ _074_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__and4_1
X_217_ net28 net27 div_q\[2\] VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__or3_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_148_ _111_ _115_ net25 _110_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__a2bb2o_1
Xoutput18 net18 VGND VGND VPWR VPWR cycl_count_o[3] sky130_fd_sc_hd__buf_2
XFILLER_7_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout31 net12 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_4
X_181_ net5 div_q\[3\] VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_13_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_250_ _078_ _079_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__a21oi_4
X_164_ net24 VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__inv_2
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_302_ net33 _021_ net30 VGND VGND VPWR VPWR div_q\[5\] sky130_fd_sc_hd__dfrtp_1
X_233_ _057_ _058_ _076_ _077_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__o211a_1
XFILLER_10_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_216_ net22 _060_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__xnor2_1
X_147_ net26 _114_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__nand2_1
Xoutput19 net19 VGND VGND VPWR VPWR cycl_count_o[4] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_15_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_18_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout32 net12 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_13_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_180_ net2 _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_3_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_163_ _129_ _130_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__nand2b_2
X_232_ net21 _059_ _075_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand3_1
X_301_ net33 _020_ net30 VGND VGND VPWR VPWR div_q\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_1_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_146_ net28 net27 div_q\[2\] div_q\[3\] VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__and4_1
X_215_ div_q\[4\] div_q\[5\] div_q\[6\] _054_ div_q\[7\] VGND VGND VPWR VPWR _060_
+ sky130_fd_sc_hd__o41a_1
XFILLER_21_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout33 net34 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XFILLER_1_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_162_ clk_gate_state_q\[1\] clk_gate_state_q\[0\] VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__and2b_1
X_300_ net33 _019_ net30 VGND VGND VPWR VPWR div_q\[3\] sky130_fd_sc_hd__dfrtp_4
X_231_ _059_ _075_ net21 VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__a21o_1
XFILLER_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 clk_i VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_145_ net28 net27 div_q\[2\] VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__and3_1
X_214_ net26 net25 div_q\[6\] _054_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__or4_1
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout34 net1 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_161_ clk_div_bypass_en_q gate_is_open_q VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__and2b_1
X_230_ net26 net25 _054_ div_q\[6\] VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__o31ai_1
XTAP_TAPCELL_ROW_19_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 div_i[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_19_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_144_ net28 net27 VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__nand2_1
X_213_ _055_ _056_ net20 VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__a21boi_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout24 _131_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout35 net1 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_1
X_160_ div_q\[3\] net17 VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ net34 _008_ net31 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dfrtp_1
Xinput3 div_i[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_10_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_143_ div_q\[6\] net20 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__xor2_1
X_212_ net20 _055_ _056_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__and3b_1
XFILLER_21_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout25 div_q\[5\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
X_288_ net34 _007_ net31 VGND VGND VPWR VPWR even_clk sky130_fd_sc_hd__dfrtp_1
Xinput4 div_i[2] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_10_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_142_ net34 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__inv_2
X_211_ net26 _054_ net25 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_10_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout26 div_q\[4\] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_2
X_287_ _003_ _006_ net31 VGND VGND VPWR VPWR i_odd_clk_xor.clk1_i sky130_fd_sc_hd__dfrtp_1
Xinput5 div_i[3] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_141_ net19 VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__inv_2
X_210_ net26 net25 _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__or3_1
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout27 div_q\[1\] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
X_286_ _002_ i_clk_gate.en_i net31 VGND VGND VPWR VPWR gate_is_open_q sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 div_i[4] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_140_ div_q\[7\] VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_269_ net21 _102_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__or2_1
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout28 div_q\[0\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_2
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_285_ net33 _005_ net30 VGND VGND VPWR VPWR clk_gate_state_q\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 div_i[5] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
X_199_ i_odd_clk_xor.clk1_i i_clk_mux.clk_sel_i VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nand2_1
X_268_ net21 _102_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand2_1
XFILLER_21_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput10 div_valid_i VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_22_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout29 net15 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_2
X_284_ net33 _004_ net30 VGND VGND VPWR VPWR clk_gate_state_q\[0\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_17_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput8 div_i[6] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_8
XPHY_EDGE_ROW_2_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_198_ clk_div_bypass_en_q net13 VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__nor2_1
X_267_ _093_ _103_ _104_ _091_ net20 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a32o_1
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 en_i VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_21_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_283_ i_clk_mux.clk_sel_i net24 _108_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__a21o_1
Xinput9 div_i[7] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_8
X_197_ _049_ _030_ net10 _132_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__a31o_1
XFILLER_18_104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_266_ net19 _097_ net20 VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_249_ clk_div_bypass_en_q _132_ _091_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__or3_1
Xinput12 rst_ni VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_282_ _032_ clk_div_bypass_en_q _131_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__mux2_1
XFILLER_18_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_196_ _048_ _047_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nor2_2
X_265_ _102_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__inv_2
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput13 test_mode_en_i VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_179_ net6 net36 net37 _031_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nor4_4
X_248_ clk_gate_state_q\[1\] _133_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_22_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_281_ net9 div_q\[7\] _131_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__mux2_1
XFILLER_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_195_ net28 _033_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__xnor2_2
X_264_ net19 net20 _097_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_6_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_247_ even_clk _090_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__xnor2_1
X_178_ net3 net5 net4 net7 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__or4_4
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ net38 div_q\[6\] net24 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__mux2_1
XFILLER_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_263_ _093_ _100_ _101_ _091_ net19 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a32o_1
X_194_ _046_ _040_ _041_ _039_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__or4_4
X_177_ clk_gate_state_q\[0\] clk_gate_state_q\[1\] VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nor2_1
X_246_ _086_ _089_ net22 _136_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__a211o_1
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_229_ div_q\[7\] _059_ _066_ _067_ _070_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__o2111a_1
XFILLER_17_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_193_ _043_ _042_ _044_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__a22o_1
X_262_ net19 _097_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__or2_1
X_176_ i_odd_clk_xor.clk1_i _029_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__xor2_1
X_245_ net17 net18 _087_ _088_ VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__or4_1
XFILLER_22_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_228_ net17 _069_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__xnor2_1
X_159_ _109_ net21 net22 VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__o21ai_1
XFILLER_17_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_261_ net19 _097_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__nand2_1
X_192_ net7 net25 VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nand2_1
XFILLER_11_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_244_ net19 net20 net21 VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__or3_1
X_175_ _119_ _123_ _135_ _028_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__and4_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_158_ _112_ _125_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__xor2_1
X_227_ _110_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__xnor2_1
XFILLER_3_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_260_ _093_ _098_ _099_ _091_ net18 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__a32o_1
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_191_ net7 net25 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__or2_1
XFILLER_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_243_ net29 net16 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__or2_1
X_174_ _113_ _128_ _026_ _027_ _126_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__o2111a_1
XFILLER_20_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_157_ div_q\[2\] net16 VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__xor2_1
X_226_ net26 _054_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__xor2_1
XFILLER_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_209_ net28 net27 div_q\[2\] div_q\[3\] VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__or4_2
XPHY_EDGE_ROW_13_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_190_ net9 div_q\[7\] VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_1_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_173_ _114_ _124_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__xnor2_1
X_242_ _124_ _125_ _081_ _085_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__or4_1
XFILLER_20_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_225_ net16 _137_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__xor2_1
XFILLER_8_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_156_ net26 net18 VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__xor2_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_208_ _129_ _130_ _030_ _053_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__a22o_1
XFILLER_15_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_172_ i_clk_mux.clk_sel_i _127_ _138_ _139_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and4_1
X_241_ _117_ _084_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__nand2_1
XFILLER_22_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_224_ _062_ _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nand2_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_155_ _122_ _121_ _120_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__mux2_1
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_207_ net13 i_clk_gate.en_i VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_171_ _113_ _128_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__nand2_1
X_240_ div_q\[5\] _110_ _082_ _083_ i_clk_mux.clk_sel_i VGND VGND VPWR VPWR _084_
+ sky130_fd_sc_hd__a221oi_1
Xrebuffer1 net9 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_223_ net28 net27 div_q\[2\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__o21ai_1
X_154_ div_q\[7\] net21 VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__xnor2_1
X_206_ i_clk_gate.clk_en _002_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__and2_1
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_170_ net29 _137_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__xnor2_1
X_299_ net33 _018_ net30 VGND VGND VPWR VPWR div_q\[2\] sky130_fd_sc_hd__dfrtp_4
Xrebuffer2 net8 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_222_ _062_ _063_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand2_1
X_153_ _109_ net21 net22 VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__a21o_1
XFILLER_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ _053_ _030_ VGND VGND VPWR VPWR gate_en_d sky130_fd_sc_hd__and2b_1
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_62 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_298_ net33 _017_ net30 VGND VGND VPWR VPWR div_q\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_9_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer3 net8 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlymetal6s4s_1
XTAP_TAPCELL_ROW_12_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_221_ _062_ _063_ _064_ _065_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__o211a_1
X_152_ net26 net25 div_q\[6\] _114_ VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__and4_1
X_204_ _047_ _048_ net10 VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__o21a_1
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_2_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_297_ net33 _016_ net30 VGND VGND VPWR VPWR div_q\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_220_ net28 net29 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__or2_1
XFILLER_12_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_151_ _117_ _118_ _116_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__mux2_1
X_203_ net11 gate_en_q VGND VGND VPWR VPWR i_clk_gate.en_i sky130_fd_sc_hd__and2_1
XFILLER_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_296_ net35 _015_ net32 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_4
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_150_ _115_ _117_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_279_ net7 net25 _131_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__mux2_1
X_202_ _002_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__inv_2
XFILLER_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_295_ net35 _014_ net32 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_4
XTAP_TAPCELL_ROW_8_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_278_ net6 net26 net24 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__mux2_1
X_201_ net34 _052_ _050_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__mux2_1
XFILLER_9_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

