* NGSPICE file created from freq_psc.ext - technology: sky130A
.subckt freq_psc VGND VPWR clk out psc[0] psc[1] psc[2] psc[3] psc[4] psc[5] psc[6] psc[7] psc[8] psc[9]
+psc[10] psc[11] psc[12] psc[13] psc[14] psc[15] rst
X_200_ psc_cnt\[12\] _076_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__or2_1
X_131_ _097_ _099_ _096_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_5_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_114_ net6 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__inv_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ net5 _085_ _086_ net4 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_8_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_113_ psc_cnt\[15\] VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_189_ psc_cnt\[8\] _069_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__or2_1
XFILLER_9_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_188_ _069_ net20 _067_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__and3b_1
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_92 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_187_ _089_ _065_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nor2_1
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload0 clknet_1_1__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_2
XFILLER_1_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_239_ clknet_1_0__leaf_clk _004_ _029_ VGND VGND VPWR VPWR psc_cnt\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_186_ psc_cnt\[7\] psc_cnt\[6\] VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__and2_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_169_ psc_cnt\[1\] psc_cnt\[0\] psc_cnt\[2\] VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a21o_1
X_238_ clknet_1_0__leaf_clk _003_ _028_ VGND VGND VPWR VPWR psc_cnt\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_185_ _089_ _065_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand2_1
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_168_ net23 _054_ _055_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__and3_1
X_237_ clknet_1_1__leaf_clk _002_ _027_ VGND VGND VPWR VPWR psc_cnt\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_13_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_184_ net20 _065_ _066_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and3_1
X_167_ psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__nand2_1
X_236_ clknet_1_1__leaf_clk _001_ _026_ VGND VGND VPWR VPWR psc_cnt\[10\] sky130_fd_sc_hd__dfrtp_1
X_219_ net22 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_11_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_183_ psc_cnt\[6\] _064_ VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_9_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_235_ clknet_1_1__leaf_clk _015_ _025_ VGND VGND VPWR VPWR psc_cnt\[9\] sky130_fd_sc_hd__dfrtp_1
X_166_ psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__or2_1
X_149_ psc_cnt\[4\] _091_ _092_ psc_cnt\[3\] _038_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__o221a_1
X_218_ net22 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ psc_cnt\[6\] _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nand2_1
XFILLER_13_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_165_ psc_cnt\[0\] net19 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and2b_1
X_234_ clknet_1_1__leaf_clk _014_ _024_ VGND VGND VPWR VPWR psc_cnt\[8\] sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_7_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_148_ psc_cnt\[7\] net14 VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__nand2b_1
X_217_ net22 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
XFILLER_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_181_ _064_ net20 _062_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__and3b_1
Xfanout20 _053_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_6
XFILLER_13_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_233_ clknet_1_1__leaf_clk _013_ _023_ VGND VGND VPWR VPWR psc_cnt\[7\] sky130_fd_sc_hd__dfrtp_1
X_164_ net26 net23 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_147_ _035_ _036_ _034_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21o_1
X_216_ net22 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout21 net17 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
X_180_ _059_ _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__and2_1
XFILLER_13_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_232_ clknet_1_1__leaf_clk _012_ _022_ VGND VGND VPWR VPWR psc_cnt\[6\] sky130_fd_sc_hd__dfrtp_1
X_163_ _052_ _049_ _051_ _101_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__o211a_4
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_146_ _093_ psc_cnt\[2\] _094_ psc_cnt\[1\] VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__o22a_1
X_215_ net22 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__inv_2
XFILLER_7_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_129_ net24 net7 VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__and2b_1
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout22 net17 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_231_ clknet_1_1__leaf_clk _011_ _021_ VGND VGND VPWR VPWR psc_cnt\[5\] sky130_fd_sc_hd__dfrtp_1
X_162_ _050_ _103_ _107_ _110_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__or4b_4
Xinput1 psc[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_145_ _094_ psc_cnt\[1\] _095_ psc_cnt\[0\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__a211o_1
X_214_ net22 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__inv_2
X_128_ _084_ psc_cnt\[14\] net5 _085_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_230_ clknet_1_0__leaf_clk _010_ _020_ VGND VGND VPWR VPWR psc_cnt\[4\] sky130_fd_sc_hd__dfrtp_1
X_161_ _103_ _112_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__or2_1
XFILLER_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 psc[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_144_ _092_ psc_cnt\[3\] _093_ psc_cnt\[2\] VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ net21 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_127_ net7 _083_ _084_ psc_cnt\[14\] VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__a2bb2o_4
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_14_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_160_ _088_ net15 _109_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a21o_1
Xinput3 psc[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_212_ net21 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_6_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_143_ _107_ _109_ _110_ _111_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__o31a_1
X_126_ net21 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 psc[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_211_ net21 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__inv_2
XFILLER_10_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_142_ _104_ _105_ _106_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__a21bo_1
X_125_ net1 VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__inv_2
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput5 psc[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_210_ net21 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__inv_2
X_141_ net16 _087_ _088_ net15 VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__o22a_1
X_124_ net8 VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__inv_2
XFILLER_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput6 psc[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_140_ _104_ _105_ _106_ _108_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__nand4_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ net9 VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__inv_2
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 psc[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_199_ _076_ net20 _075_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__and3b_1
X_122_ net10 VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__inv_2
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput10 psc[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 psc[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_198_ psc_cnt\[11\] psc_cnt\[10\] psc_cnt\[9\] _071_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__and4_1
XFILLER_2_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_121_ net11 VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__inv_2
Xinput11 psc[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout19 _053_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_6
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 psc[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_197_ psc_cnt\[10\] psc_cnt\[9\] _071_ psc_cnt\[11\] VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__a31o_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ psc_cnt\[6\] VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__inv_2
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput12 psc[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_196_ net20 _074_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__and2_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 psc[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_179_ psc_cnt\[5\] psc_cnt\[4\] VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_10_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_13_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_195_ psc_cnt\[10\] _072_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__xnor2_1
Xinput14 psc[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
X_178_ psc_cnt\[4\] _059_ psc_cnt\[5\] VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__a21o_1
XFILLER_8_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ _073_ net20 _072_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_11_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput15 psc[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_177_ net19 _060_ _061_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__and3_1
XFILLER_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_229_ clknet_1_0__leaf_clk _009_ _019_ VGND VGND VPWR VPWR psc_cnt\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 net18 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_193_ psc_cnt\[9\] _071_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__nor2_1
Xinput16 psc[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_176_ psc_cnt\[4\] _059_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_159_ _037_ _046_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__a21oi_1
X_228_ clknet_1_0__leaf_clk _008_ _018_ VGND VGND VPWR VPWR psc_cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_17_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclone1 _053_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_6
XFILLER_17_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold5 _083_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_17_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_192_ psc_cnt\[9\] _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nand2_1
XFILLER_2_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 rst VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
X_175_ psc_cnt\[4\] _059_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_5_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_158_ _043_ _047_ _038_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__a21boi_1
X_227_ clknet_1_0__leaf_clk _007_ _017_ VGND VGND VPWR VPWR psc_cnt\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ _071_ net20 _070_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__and3b_1
X_174_ _059_ net19 _058_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__and3b_1
X_157_ net13 _090_ _040_ _041_ _044_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__a221o_1
X_226_ clknet_1_0__leaf_clk _000_ _016_ VGND VGND VPWR VPWR psc_cnt\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_209_ net27 _082_ net23 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__a21boi_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ psc_cnt\[8\] _059_ _063_ _068_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__and4_1
X_173_ psc_cnt\[3\] psc_cnt\[2\] psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _059_
+ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_7_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_242_ clknet_1_0__leaf_clk _033_ _032_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_3_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_156_ _039_ _042_ _043_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__and4_1
X_225_ net21 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_208_ net19 _081_ _082_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__and3_1
X_139_ psc_cnt\[10\] net2 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_172_ psc_cnt\[2\] psc_cnt\[1\] psc_cnt\[0\] psc_cnt\[3\] VGND VGND VPWR VPWR _058_
+ sky130_fd_sc_hd__a31o_1
X_241_ clknet_1_0__leaf_clk _006_ _031_ VGND VGND VPWR VPWR psc_cnt\[15\] sky130_fd_sc_hd__dfrtp_1
X_155_ net13 _090_ _044_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a21oi_1
X_224_ net21 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_9_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_207_ net25 _079_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__nand2_1
X_138_ net16 _087_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__and2_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_171_ net23 _056_ _057_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__and3_1
X_240_ clknet_1_0__leaf_clk _005_ _030_ VGND VGND VPWR VPWR psc_cnt\[14\] sky130_fd_sc_hd__dfrtp_1
X_223_ net21 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
X_154_ psc_cnt\[5\] net12 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and2b_1
XFILLER_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_206_ psc_cnt\[14\] _079_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__or2_1
X_137_ psc_cnt\[11\] net3 VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ psc_cnt\[2\] psc_cnt\[1\] psc_cnt\[0\] VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nand3_1
Xrebuffer2 psc_cnt\[15\] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
X_153_ net14 _089_ net13 _090_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_8_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ net21 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
XFILLER_12_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_205_ net23 _080_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and2_1
X_136_ net3 psc_cnt\[11\] VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_119_ psc_cnt\[7\] VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrebuffer3 psc_cnt\[14\] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_152_ _040_ _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2_1
X_221_ net21 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
X_204_ _085_ _078_ _079_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_135_ net2 psc_cnt\[10\] VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__nand2b_1
X_118_ psc_cnt\[8\] VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__inv_2
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_151_ net11 psc_cnt\[4\] VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nand2b_1
X_220_ net22 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__inv_2
XFILLER_17_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_203_ psc_cnt\[13\] psc_cnt\[12\] _076_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__and3_1
X_134_ _097_ _096_ _099_ _102_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__or4bb_4
X_117_ psc_cnt\[9\] VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__inv_2
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_1_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_150_ net12 psc_cnt\[5\] VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2b_1
XFILLER_6_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_4_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ net19 _077_ _078_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and3_1
X_133_ _086_ net4 _098_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__a21oi_1
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_116_ psc_cnt\[12\] VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_201_ psc_cnt\[12\] _076_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__nand2_1
X_132_ _098_ _100_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__or2_1
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_115_ psc_cnt\[13\] VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__inv_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
.ends

