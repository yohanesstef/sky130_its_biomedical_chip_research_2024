magic
tech sky130A
magscale 1 2
timestamp 1730101540
<< viali >>
rect 9045 13957 9079 13991
rect 5273 13889 5307 13923
rect 6101 13889 6135 13923
rect 6561 13889 6595 13923
rect 7205 13889 7239 13923
rect 7941 13889 7975 13923
rect 9321 13889 9355 13923
rect 9873 13889 9907 13923
rect 8493 13821 8527 13855
rect 10149 13821 10183 13855
rect 5457 13753 5491 13787
rect 9229 13753 9263 13787
rect 5917 13685 5951 13719
rect 6745 13685 6779 13719
rect 7389 13685 7423 13719
rect 9505 13685 9539 13719
rect 6653 13481 6687 13515
rect 8401 13481 8435 13515
rect 5641 13413 5675 13447
rect 7849 13413 7883 13447
rect 6101 13345 6135 13379
rect 7757 13345 7791 13379
rect 7978 13345 8012 13379
rect 8493 13345 8527 13379
rect 9689 13345 9723 13379
rect 3985 13277 4019 13311
rect 4077 13277 4111 13311
rect 4169 13277 4203 13311
rect 6009 13277 6043 13311
rect 6561 13277 6595 13311
rect 6653 13277 6687 13311
rect 7113 13277 7147 13311
rect 8579 13277 8613 13311
rect 9597 13277 9631 13311
rect 7297 13209 7331 13243
rect 8125 13209 8159 13243
rect 4353 13141 4387 13175
rect 6285 13141 6319 13175
rect 6929 13141 6963 13175
rect 7481 13141 7515 13175
rect 8217 13141 8251 13175
rect 9965 13141 9999 13175
rect 4629 12937 4663 12971
rect 7205 12937 7239 12971
rect 8309 12937 8343 12971
rect 9965 12937 9999 12971
rect 7389 12869 7423 12903
rect 7573 12869 7607 12903
rect 8493 12869 8527 12903
rect 10149 12869 10183 12903
rect 3801 12801 3835 12835
rect 4169 12801 4203 12835
rect 4261 12801 4295 12835
rect 4445 12801 4479 12835
rect 4721 12801 4755 12835
rect 5089 12801 5123 12835
rect 5549 12801 5583 12835
rect 6193 12801 6227 12835
rect 6653 12801 6687 12835
rect 6929 12801 6963 12835
rect 7021 12801 7055 12835
rect 7297 12801 7331 12835
rect 7665 12801 7699 12835
rect 7757 12801 7791 12835
rect 7941 12801 7975 12835
rect 8033 12801 8067 12835
rect 8125 12801 8159 12835
rect 8677 12801 8711 12835
rect 8769 12801 8803 12835
rect 9045 12801 9079 12835
rect 9137 12801 9171 12835
rect 9413 12801 9447 12835
rect 9873 12801 9907 12835
rect 10057 12801 10091 12835
rect 10701 12801 10735 12835
rect 10885 12801 10919 12835
rect 3893 12733 3927 12767
rect 4997 12733 5031 12767
rect 5411 12733 5445 12767
rect 6837 12733 6871 12767
rect 8953 12733 8987 12767
rect 4353 12665 4387 12699
rect 4813 12665 4847 12699
rect 6469 12665 6503 12699
rect 7389 12665 7423 12699
rect 10517 12665 10551 12699
rect 10793 12665 10827 12699
rect 3525 12597 3559 12631
rect 4905 12597 4939 12631
rect 5181 12597 5215 12631
rect 5273 12597 5307 12631
rect 5733 12597 5767 12631
rect 6745 12597 6779 12631
rect 7021 12597 7055 12631
rect 9229 12597 9263 12631
rect 9505 12597 9539 12631
rect 10609 12597 10643 12631
rect 3065 12393 3099 12427
rect 3525 12393 3559 12427
rect 4077 12393 4111 12427
rect 5917 12393 5951 12427
rect 6929 12393 6963 12427
rect 11345 12393 11379 12427
rect 6028 12325 6062 12359
rect 8309 12325 8343 12359
rect 10609 12325 10643 12359
rect 4537 12257 4571 12291
rect 5825 12257 5859 12291
rect 7849 12257 7883 12291
rect 10793 12257 10827 12291
rect 3249 12189 3283 12223
rect 3341 12189 3375 12223
rect 3617 12189 3651 12223
rect 4261 12189 4295 12223
rect 4445 12189 4479 12223
rect 4629 12191 4663 12225
rect 4813 12189 4847 12223
rect 6193 12189 6227 12223
rect 6745 12189 6779 12223
rect 6929 12189 6963 12223
rect 7941 12189 7975 12223
rect 8401 12189 8435 12223
rect 9137 12189 9171 12223
rect 9229 12189 9263 12223
rect 9505 12189 9539 12223
rect 9781 12189 9815 12223
rect 10057 12189 10091 12223
rect 10241 12189 10275 12223
rect 10425 12189 10459 12223
rect 10701 12189 10735 12223
rect 10977 12189 11011 12223
rect 11069 12189 11103 12223
rect 11529 12189 11563 12223
rect 11805 12189 11839 12223
rect 9321 12121 9355 12155
rect 10333 12121 10367 12155
rect 5549 12053 5583 12087
rect 8493 12053 8527 12087
rect 8953 12053 8987 12087
rect 9689 12053 9723 12087
rect 11253 12053 11287 12087
rect 11713 12053 11747 12087
rect 6469 11849 6503 11883
rect 11529 11849 11563 11883
rect 12341 11849 12375 11883
rect 12541 11781 12575 11815
rect 3249 11713 3283 11747
rect 3985 11713 4019 11747
rect 4077 11713 4111 11747
rect 4169 11713 4203 11747
rect 4353 11713 4387 11747
rect 4905 11713 4939 11747
rect 5089 11713 5123 11747
rect 5181 11713 5215 11747
rect 5273 11713 5307 11747
rect 5391 11713 5425 11747
rect 5825 11713 5859 11747
rect 6009 11713 6043 11747
rect 6377 11713 6411 11747
rect 7941 11713 7975 11747
rect 8217 11713 8251 11747
rect 8309 11713 8343 11747
rect 9229 11713 9263 11747
rect 9321 11713 9355 11747
rect 9597 11713 9631 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 11897 11713 11931 11747
rect 12081 11713 12115 11747
rect 3341 11645 3375 11679
rect 3433 11645 3467 11679
rect 3709 11645 3743 11679
rect 5549 11645 5583 11679
rect 8033 11645 8067 11679
rect 9505 11645 9539 11679
rect 3617 11577 3651 11611
rect 3433 11509 3467 11543
rect 5641 11509 5675 11543
rect 8493 11509 8527 11543
rect 9045 11509 9079 11543
rect 12173 11509 12207 11543
rect 12357 11509 12391 11543
rect 3893 11305 3927 11339
rect 4445 11305 4479 11339
rect 11529 11305 11563 11339
rect 8493 11169 8527 11203
rect 11345 11169 11379 11203
rect 4077 11101 4111 11135
rect 4261 11101 4295 11135
rect 4353 11101 4387 11135
rect 4629 11101 4663 11135
rect 4997 11101 5031 11135
rect 5549 11101 5583 11135
rect 5825 11101 5859 11135
rect 8309 11101 8343 11135
rect 9413 11101 9447 11135
rect 9597 11101 9631 11135
rect 11805 11101 11839 11135
rect 12173 11101 12207 11135
rect 12909 11101 12943 11135
rect 4721 11033 4755 11067
rect 4813 11033 4847 11067
rect 12449 11033 12483 11067
rect 5457 10965 5491 10999
rect 5917 10965 5951 10999
rect 8125 10965 8159 10999
rect 9505 10965 9539 10999
rect 11713 10965 11747 10999
rect 11989 10965 12023 10999
rect 12357 10761 12391 10795
rect 6009 10693 6043 10727
rect 8217 10693 8251 10727
rect 11529 10693 11563 10727
rect 12265 10693 12299 10727
rect 5549 10625 5583 10659
rect 5641 10625 5675 10659
rect 6929 10625 6963 10659
rect 8033 10625 8067 10659
rect 8309 10625 8343 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 9321 10625 9355 10659
rect 9689 10625 9723 10659
rect 12541 10625 12575 10659
rect 12725 10625 12759 10659
rect 12817 10625 12851 10659
rect 1501 10557 1535 10591
rect 3249 10557 3283 10591
rect 3525 10557 3559 10591
rect 5917 10557 5951 10591
rect 6745 10557 6779 10591
rect 6837 10557 6871 10591
rect 8585 10557 8619 10591
rect 8769 10557 8803 10591
rect 8861 10557 8895 10591
rect 9413 10557 9447 10591
rect 10333 10557 10367 10591
rect 11897 10557 11931 10591
rect 6561 10489 6595 10523
rect 9229 10489 9263 10523
rect 10057 10489 10091 10523
rect 11989 10489 12023 10523
rect 5365 10421 5399 10455
rect 6745 10421 6779 10455
rect 7849 10421 7883 10455
rect 9597 10421 9631 10455
rect 9873 10421 9907 10455
rect 12127 10421 12161 10455
rect 3525 10217 3559 10251
rect 3893 10217 3927 10251
rect 9505 10217 9539 10251
rect 10333 10217 10367 10251
rect 10885 10217 10919 10251
rect 12449 10217 12483 10251
rect 12817 10217 12851 10251
rect 7021 10149 7055 10183
rect 8677 10149 8711 10183
rect 8953 10149 8987 10183
rect 10425 10149 10459 10183
rect 11529 10149 11563 10183
rect 11713 10149 11747 10183
rect 1777 10081 1811 10115
rect 4261 10081 4295 10115
rect 5365 10081 5399 10115
rect 9229 10081 9263 10115
rect 12541 10081 12575 10115
rect 1501 10013 1535 10047
rect 1685 10013 1719 10047
rect 3985 10013 4019 10047
rect 4169 10013 4203 10047
rect 4445 10013 4479 10047
rect 4537 10013 4571 10047
rect 4813 10013 4847 10047
rect 5273 10013 5307 10047
rect 5641 10013 5675 10047
rect 5733 10013 5767 10047
rect 6285 10013 6319 10047
rect 6469 10013 6503 10047
rect 6561 10013 6595 10047
rect 6653 10013 6687 10047
rect 7021 10013 7055 10047
rect 7297 10013 7331 10047
rect 7481 10013 7515 10047
rect 8125 10013 8159 10047
rect 8217 10013 8251 10047
rect 9137 10013 9171 10047
rect 9689 10013 9723 10047
rect 9782 10013 9816 10047
rect 10195 10013 10229 10047
rect 10609 10013 10643 10047
rect 10701 10013 10735 10047
rect 10977 10013 11011 10047
rect 11069 10013 11103 10047
rect 11851 10013 11885 10047
rect 12209 10013 12243 10047
rect 12357 10013 12391 10047
rect 12449 10013 12483 10047
rect 2053 9945 2087 9979
rect 4997 9945 5031 9979
rect 7941 9945 7975 9979
rect 8677 9945 8711 9979
rect 9597 9945 9631 9979
rect 9965 9945 9999 9979
rect 10057 9945 10091 9979
rect 11989 9945 12023 9979
rect 12081 9945 12115 9979
rect 1685 9877 1719 9911
rect 4721 9877 4755 9911
rect 6929 9877 6963 9911
rect 7205 9877 7239 9911
rect 7573 9877 7607 9911
rect 2053 9673 2087 9707
rect 3617 9673 3651 9707
rect 4905 9673 4939 9707
rect 7205 9673 7239 9707
rect 9321 9673 9355 9707
rect 10517 9673 10551 9707
rect 12081 9673 12115 9707
rect 1593 9605 1627 9639
rect 1777 9605 1811 9639
rect 2237 9605 2271 9639
rect 3769 9605 3803 9639
rect 3985 9605 4019 9639
rect 4169 9605 4203 9639
rect 5917 9605 5951 9639
rect 10241 9605 10275 9639
rect 11161 9605 11195 9639
rect 1961 9537 1995 9571
rect 2881 9537 2915 9571
rect 3065 9537 3099 9571
rect 3341 9537 3375 9571
rect 4261 9537 4295 9571
rect 4629 9537 4663 9571
rect 4721 9537 4755 9571
rect 5365 9537 5399 9571
rect 5549 9537 5583 9571
rect 5825 9537 5859 9571
rect 6009 9537 6043 9571
rect 6101 9537 6135 9571
rect 6377 9537 6411 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 7205 9537 7239 9571
rect 7389 9537 7423 9571
rect 9229 9537 9263 9571
rect 9321 9537 9355 9571
rect 9505 9537 9539 9571
rect 10701 9537 10735 9571
rect 10793 9537 10827 9571
rect 11069 9537 11103 9571
rect 11621 9537 11655 9571
rect 11989 9537 12023 9571
rect 12265 9537 12299 9571
rect 12449 9537 12483 9571
rect 12725 9537 12759 9571
rect 12817 9537 12851 9571
rect 2605 9469 2639 9503
rect 3157 9469 3191 9503
rect 3525 9469 3559 9503
rect 5641 9469 5675 9503
rect 8677 9469 8711 9503
rect 9781 9469 9815 9503
rect 11713 9469 11747 9503
rect 12541 9469 12575 9503
rect 5365 9401 5399 9435
rect 8769 9401 8803 9435
rect 9965 9401 9999 9435
rect 11805 9401 11839 9435
rect 2237 9333 2271 9367
rect 2697 9333 2731 9367
rect 3801 9333 3835 9367
rect 7021 9333 7055 9367
rect 8401 9333 8435 9367
rect 8861 9333 8895 9367
rect 11897 9333 11931 9367
rect 12633 9333 12667 9367
rect 3341 9129 3375 9163
rect 9413 9129 9447 9163
rect 11345 9129 11379 9163
rect 12541 9129 12575 9163
rect 12817 9129 12851 9163
rect 6377 9061 6411 9095
rect 2789 8993 2823 9027
rect 2881 8993 2915 9027
rect 2697 8925 2731 8959
rect 2973 8925 3007 8959
rect 4813 8925 4847 8959
rect 6285 8925 6319 8959
rect 6561 8925 6595 8959
rect 6653 8925 6687 8959
rect 9229 8925 9263 8959
rect 9413 8925 9447 8959
rect 11253 8925 11287 8959
rect 12725 8925 12759 8959
rect 13001 8925 13035 8959
rect 3309 8857 3343 8891
rect 3525 8857 3559 8891
rect 4997 8857 5031 8891
rect 2513 8789 2547 8823
rect 3157 8789 3191 8823
rect 4629 8789 4663 8823
rect 6837 8789 6871 8823
rect 3617 8585 3651 8619
rect 2145 8517 2179 8551
rect 5917 8517 5951 8551
rect 12357 8517 12391 8551
rect 6009 8449 6043 8483
rect 10701 8449 10735 8483
rect 12633 8449 12667 8483
rect 12725 8449 12759 8483
rect 1869 8381 1903 8415
rect 3985 8381 4019 8415
rect 4261 8381 4295 8415
rect 5733 8381 5767 8415
rect 10609 8381 10643 8415
rect 11161 8381 11195 8415
rect 12817 8313 12851 8347
rect 2237 8041 2271 8075
rect 2421 8041 2455 8075
rect 2973 8041 3007 8075
rect 7389 8041 7423 8075
rect 8033 8041 8067 8075
rect 8677 8041 8711 8075
rect 10517 8041 10551 8075
rect 12541 8041 12575 8075
rect 4261 7973 4295 8007
rect 7665 7973 7699 8007
rect 8953 7973 8987 8007
rect 5641 7905 5675 7939
rect 9505 7905 9539 7939
rect 11069 7905 11103 7939
rect 1869 7837 1903 7871
rect 2881 7837 2915 7871
rect 3525 7837 3559 7871
rect 8493 7837 8527 7871
rect 10793 7837 10827 7871
rect 12725 7837 12759 7871
rect 5549 7769 5583 7803
rect 5917 7769 5951 7803
rect 8309 7769 8343 7803
rect 9321 7769 9355 7803
rect 10333 7769 10367 7803
rect 12817 7769 12851 7803
rect 2237 7701 2271 7735
rect 8033 7701 8067 7735
rect 8217 7701 8251 7735
rect 9137 7701 9171 7735
rect 9229 7701 9263 7735
rect 10533 7701 10567 7735
rect 10701 7701 10735 7735
rect 4445 7497 4479 7531
rect 4705 7497 4739 7531
rect 6745 7497 6779 7531
rect 9413 7497 9447 7531
rect 11069 7497 11103 7531
rect 4261 7429 4295 7463
rect 4905 7429 4939 7463
rect 6193 7429 6227 7463
rect 7941 7429 7975 7463
rect 9597 7429 9631 7463
rect 11529 7429 11563 7463
rect 11713 7429 11747 7463
rect 5641 7361 5675 7395
rect 6009 7361 6043 7395
rect 6653 7361 6687 7395
rect 7665 7361 7699 7395
rect 9689 7361 9723 7395
rect 11069 7361 11103 7395
rect 11263 7361 11297 7395
rect 11897 7361 11931 7395
rect 5365 7293 5399 7327
rect 12541 7293 12575 7327
rect 3893 7225 3927 7259
rect 4537 7225 4571 7259
rect 4261 7157 4295 7191
rect 4721 7157 4755 7191
rect 5825 7157 5859 7191
rect 12081 7157 12115 7191
rect 5365 6953 5399 6987
rect 5549 6953 5583 6987
rect 7757 6953 7791 6987
rect 8309 6953 8343 6987
rect 8493 6953 8527 6987
rect 11326 6953 11360 6987
rect 12817 6953 12851 6987
rect 6101 6885 6135 6919
rect 4813 6817 4847 6851
rect 8953 6817 8987 6851
rect 11069 6817 11103 6851
rect 1409 6749 1443 6783
rect 2145 6749 2179 6783
rect 2881 6749 2915 6783
rect 4721 6749 4755 6783
rect 4997 6749 5031 6783
rect 5641 6749 5675 6783
rect 5825 6749 5859 6783
rect 6009 6749 6043 6783
rect 6285 6749 6319 6783
rect 6469 6749 6503 6783
rect 2329 6681 2363 6715
rect 8477 6681 8511 6715
rect 8677 6681 8711 6715
rect 9229 6681 9263 6715
rect 1593 6613 1627 6647
rect 2513 6613 2547 6647
rect 2973 6613 3007 6647
rect 4353 6613 4387 6647
rect 5365 6613 5399 6647
rect 10701 6613 10735 6647
rect 5733 6409 5767 6443
rect 6745 6409 6779 6443
rect 8309 6409 8343 6443
rect 9689 6409 9723 6443
rect 10399 6409 10433 6443
rect 10977 6409 11011 6443
rect 8125 6341 8159 6375
rect 8401 6341 8435 6375
rect 10609 6341 10643 6375
rect 11253 6341 11287 6375
rect 12081 6341 12115 6375
rect 1501 6273 1535 6307
rect 1593 6273 1627 6307
rect 1869 6273 1903 6307
rect 4997 6273 5031 6307
rect 5549 6273 5583 6307
rect 5641 6273 5675 6307
rect 5917 6273 5951 6307
rect 6377 6273 6411 6307
rect 6531 6273 6565 6307
rect 6837 6273 6871 6307
rect 7757 6273 7791 6307
rect 10885 6273 10919 6307
rect 11069 6273 11103 6307
rect 12633 6273 12667 6307
rect 2145 6205 2179 6239
rect 4813 6205 4847 6239
rect 5273 6205 5307 6239
rect 10701 6205 10735 6239
rect 3617 6137 3651 6171
rect 1777 6069 1811 6103
rect 5181 6069 5215 6103
rect 5365 6069 5399 6103
rect 5457 6069 5491 6103
rect 6009 6069 6043 6103
rect 6929 6069 6963 6103
rect 8125 6069 8159 6103
rect 10241 6069 10275 6103
rect 10425 6069 10459 6103
rect 2329 5865 2363 5899
rect 2513 5865 2547 5899
rect 3985 5865 4019 5899
rect 6561 5865 6595 5899
rect 7297 5865 7331 5899
rect 8677 5865 8711 5899
rect 8953 5865 8987 5899
rect 9965 5865 9999 5899
rect 10425 5865 10459 5899
rect 12633 5865 12667 5899
rect 2881 5797 2915 5831
rect 4905 5797 4939 5831
rect 7021 5797 7055 5831
rect 10793 5797 10827 5831
rect 6193 5729 6227 5763
rect 6929 5729 6963 5763
rect 10885 5729 10919 5763
rect 2145 5661 2179 5695
rect 2973 5661 3007 5695
rect 3157 5661 3191 5695
rect 4721 5661 4755 5695
rect 4997 5661 5031 5695
rect 5089 5661 5123 5695
rect 5182 5661 5216 5695
rect 5365 5661 5399 5695
rect 5593 5661 5627 5695
rect 5825 5661 5859 5695
rect 6009 5661 6043 5695
rect 6101 5661 6135 5695
rect 6377 5661 6411 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 7113 5661 7147 5695
rect 8309 5661 8343 5695
rect 8493 5661 8527 5695
rect 8585 5661 8619 5695
rect 9137 5661 9171 5695
rect 9413 5661 9447 5695
rect 9597 5661 9631 5695
rect 1777 5593 1811 5627
rect 2513 5593 2547 5627
rect 3953 5593 3987 5627
rect 4169 5593 4203 5627
rect 5457 5593 5491 5627
rect 9965 5593 9999 5627
rect 11161 5593 11195 5627
rect 3341 5525 3375 5559
rect 3801 5525 3835 5559
rect 4537 5525 4571 5559
rect 5733 5525 5767 5559
rect 8493 5525 8527 5559
rect 9321 5525 9355 5559
rect 10149 5525 10183 5559
rect 10241 5525 10275 5559
rect 10425 5525 10459 5559
rect 4813 5321 4847 5355
rect 5983 5321 6017 5355
rect 11529 5321 11563 5355
rect 12817 5321 12851 5355
rect 4261 5253 4295 5287
rect 4997 5253 5031 5287
rect 6193 5253 6227 5287
rect 8677 5253 8711 5287
rect 8893 5253 8927 5287
rect 9137 5253 9171 5287
rect 9505 5253 9539 5287
rect 11897 5253 11931 5287
rect 1869 5185 1903 5219
rect 3709 5185 3743 5219
rect 3893 5185 3927 5219
rect 3985 5185 4019 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 9321 5185 9355 5219
rect 9597 5185 9631 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 12265 5185 12299 5219
rect 12725 5185 12759 5219
rect 2145 5117 2179 5151
rect 5365 5117 5399 5151
rect 9873 5117 9907 5151
rect 11345 5117 11379 5151
rect 3893 5049 3927 5083
rect 5273 5049 5307 5083
rect 5825 5049 5859 5083
rect 3617 4981 3651 5015
rect 4261 4981 4295 5015
rect 5162 4981 5196 5015
rect 5641 4981 5675 5015
rect 6009 4981 6043 5015
rect 8861 4981 8895 5015
rect 9045 4981 9079 5015
rect 12357 4981 12391 5015
rect 2053 4777 2087 4811
rect 2237 4777 2271 4811
rect 3893 4777 3927 4811
rect 5273 4777 5307 4811
rect 6193 4777 6227 4811
rect 12265 4777 12299 4811
rect 2605 4709 2639 4743
rect 4629 4709 4663 4743
rect 6745 4709 6779 4743
rect 11897 4709 11931 4743
rect 5181 4641 5215 4675
rect 9689 4641 9723 4675
rect 3985 4573 4019 4607
rect 4813 4573 4847 4607
rect 4905 4573 4939 4607
rect 5089 4573 5123 4607
rect 6469 4573 6503 4607
rect 6561 4573 6595 4607
rect 6745 4573 6779 4607
rect 8493 4573 8527 4607
rect 8585 4573 8619 4607
rect 9413 4573 9447 4607
rect 11529 4573 11563 4607
rect 11713 4573 11747 4607
rect 12349 4573 12383 4607
rect 2237 4505 2271 4539
rect 4629 4505 4663 4539
rect 6193 4505 6227 4539
rect 7849 4505 7883 4539
rect 8033 4505 8067 4539
rect 11437 4505 11471 4539
rect 5457 4437 5491 4471
rect 6377 4437 6411 4471
rect 8217 4437 8251 4471
rect 8309 4437 8343 4471
rect 8125 4233 8159 4267
rect 8585 4165 8619 4199
rect 8801 4165 8835 4199
rect 4721 4097 4755 4131
rect 5503 4097 5537 4131
rect 6009 4097 6043 4131
rect 6193 4097 6227 4131
rect 9229 4097 9263 4131
rect 9965 4097 9999 4131
rect 10149 4097 10183 4131
rect 10333 4097 10367 4131
rect 10609 4097 10643 4131
rect 10793 4097 10827 4131
rect 10885 4097 10919 4131
rect 3893 4029 3927 4063
rect 4445 4029 4479 4063
rect 4905 4029 4939 4063
rect 4997 4029 5031 4063
rect 5365 4029 5399 4063
rect 8493 4029 8527 4063
rect 9505 4029 9539 4063
rect 5917 3961 5951 3995
rect 6101 3961 6135 3995
rect 5549 3893 5583 3927
rect 7941 3893 7975 3927
rect 8125 3893 8159 3927
rect 8769 3893 8803 3927
rect 8953 3893 8987 3927
rect 10517 3893 10551 3927
rect 5089 3689 5123 3723
rect 5825 3689 5859 3723
rect 6469 3689 6503 3723
rect 8309 3689 8343 3723
rect 9210 3689 9244 3723
rect 10701 3689 10735 3723
rect 12817 3689 12851 3723
rect 4997 3621 5031 3655
rect 4721 3553 4755 3587
rect 5273 3553 5307 3587
rect 5457 3553 5491 3587
rect 6009 3553 6043 3587
rect 8953 3553 8987 3587
rect 4629 3485 4663 3519
rect 5365 3485 5399 3519
rect 5549 3485 5583 3519
rect 6101 3485 6135 3519
rect 6561 3485 6595 3519
rect 6653 3485 6687 3519
rect 6837 3485 6871 3519
rect 6929 3485 6963 3519
rect 7113 3485 7147 3519
rect 8217 3485 8251 3519
rect 8401 3485 8435 3519
rect 8585 3485 8619 3519
rect 13001 3485 13035 3519
rect 6745 3417 6779 3451
rect 7021 3349 7055 3383
rect 8677 3349 8711 3383
rect 6101 3145 6135 3179
rect 8125 3145 8159 3179
rect 5549 3009 5583 3043
rect 6009 3009 6043 3043
rect 6193 3009 6227 3043
rect 6745 3009 6779 3043
rect 7481 3009 7515 3043
rect 7849 3009 7883 3043
rect 9873 3009 9907 3043
rect 5641 2941 5675 2975
rect 9597 2941 9631 2975
rect 6561 2873 6595 2907
rect 5825 2805 5859 2839
rect 7297 2805 7331 2839
rect 7757 2805 7791 2839
rect 5089 2601 5123 2635
rect 8217 2601 8251 2635
rect 6193 2465 6227 2499
rect 6469 2465 6503 2499
rect 5273 2397 5307 2431
rect 5917 2397 5951 2431
rect 6745 2329 6779 2363
<< metal1 >>
rect 1104 14170 13340 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 13340 14170
rect 1104 14096 13340 14118
rect 8386 13948 8392 14000
rect 8444 13988 8450 14000
rect 9033 13991 9091 13997
rect 9033 13988 9045 13991
rect 8444 13960 9045 13988
rect 8444 13948 8450 13960
rect 9033 13957 9045 13960
rect 9079 13957 9091 13991
rect 9033 13951 9091 13957
rect 5258 13880 5264 13932
rect 5316 13880 5322 13932
rect 5810 13880 5816 13932
rect 5868 13920 5874 13932
rect 6089 13923 6147 13929
rect 6089 13920 6101 13923
rect 5868 13892 6101 13920
rect 5868 13880 5874 13892
rect 6089 13889 6101 13892
rect 6135 13889 6147 13923
rect 6089 13883 6147 13889
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 6549 13923 6607 13929
rect 6549 13920 6561 13923
rect 6512 13892 6561 13920
rect 6512 13880 6518 13892
rect 6549 13889 6561 13892
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 7156 13892 7205 13920
rect 7156 13880 7162 13892
rect 7193 13889 7205 13892
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 7742 13880 7748 13932
rect 7800 13920 7806 13932
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 7800 13892 7941 13920
rect 7800 13880 7806 13892
rect 7929 13889 7941 13892
rect 7975 13889 7987 13923
rect 7929 13883 7987 13889
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 9309 13923 9367 13929
rect 9309 13920 9321 13923
rect 9180 13892 9321 13920
rect 9180 13880 9186 13892
rect 9309 13889 9321 13892
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9732 13892 9873 13920
rect 9732 13880 9738 13892
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 8294 13812 8300 13864
rect 8352 13852 8358 13864
rect 8481 13855 8539 13861
rect 8481 13852 8493 13855
rect 8352 13824 8493 13852
rect 8352 13812 8358 13824
rect 8481 13821 8493 13824
rect 8527 13852 8539 13855
rect 9398 13852 9404 13864
rect 8527 13824 9404 13852
rect 8527 13821 8539 13824
rect 8481 13815 8539 13821
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 4706 13744 4712 13796
rect 4764 13784 4770 13796
rect 5445 13787 5503 13793
rect 5445 13784 5457 13787
rect 4764 13756 5457 13784
rect 4764 13744 4770 13756
rect 5445 13753 5457 13756
rect 5491 13784 5503 13787
rect 6638 13784 6644 13796
rect 5491 13756 6644 13784
rect 5491 13753 5503 13756
rect 5445 13747 5503 13753
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 9217 13787 9275 13793
rect 9217 13753 9229 13787
rect 9263 13784 9275 13787
rect 9766 13784 9772 13796
rect 9263 13756 9772 13784
rect 9263 13753 9275 13756
rect 9217 13747 9275 13753
rect 9766 13744 9772 13756
rect 9824 13744 9830 13796
rect 9858 13744 9864 13796
rect 9916 13784 9922 13796
rect 10152 13784 10180 13815
rect 9916 13756 10180 13784
rect 9916 13744 9922 13756
rect 5902 13676 5908 13728
rect 5960 13676 5966 13728
rect 6730 13676 6736 13728
rect 6788 13676 6794 13728
rect 7190 13676 7196 13728
rect 7248 13716 7254 13728
rect 7377 13719 7435 13725
rect 7377 13716 7389 13719
rect 7248 13688 7389 13716
rect 7248 13676 7254 13688
rect 7377 13685 7389 13688
rect 7423 13685 7435 13719
rect 7377 13679 7435 13685
rect 9490 13676 9496 13728
rect 9548 13676 9554 13728
rect 1104 13626 13340 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 13340 13626
rect 1104 13552 13340 13574
rect 5810 13472 5816 13524
rect 5868 13512 5874 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 5868 13484 6653 13512
rect 5868 13472 5874 13484
rect 6641 13481 6653 13484
rect 6687 13512 6699 13515
rect 6730 13512 6736 13524
rect 6687 13484 6736 13512
rect 6687 13481 6699 13484
rect 6641 13475 6699 13481
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 8294 13512 8300 13524
rect 7760 13484 8300 13512
rect 3602 13404 3608 13456
rect 3660 13444 3666 13456
rect 5629 13447 5687 13453
rect 5629 13444 5641 13447
rect 3660 13416 5641 13444
rect 3660 13404 3666 13416
rect 5629 13413 5641 13416
rect 5675 13444 5687 13447
rect 6454 13444 6460 13456
rect 5675 13416 6460 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 6454 13404 6460 13416
rect 6512 13404 6518 13456
rect 4798 13376 4804 13388
rect 3988 13348 4804 13376
rect 3988 13317 4016 13348
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5902 13376 5908 13388
rect 5316 13348 5908 13376
rect 5316 13336 5322 13348
rect 5902 13336 5908 13348
rect 5960 13336 5966 13388
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13376 6147 13379
rect 7006 13376 7012 13388
rect 6135 13348 7012 13376
rect 6135 13345 6147 13348
rect 6089 13339 6147 13345
rect 7006 13336 7012 13348
rect 7064 13336 7070 13388
rect 7760 13385 7788 13484
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8389 13515 8447 13521
rect 8389 13481 8401 13515
rect 8435 13481 8447 13515
rect 8389 13475 8447 13481
rect 7837 13447 7895 13453
rect 7837 13413 7849 13447
rect 7883 13444 7895 13447
rect 8404 13444 8432 13475
rect 9858 13444 9864 13456
rect 7883 13416 9864 13444
rect 7883 13413 7895 13416
rect 7837 13407 7895 13413
rect 9858 13404 9864 13416
rect 9916 13404 9922 13456
rect 7745 13379 7803 13385
rect 7745 13376 7757 13379
rect 7116 13348 7757 13376
rect 3973 13311 4031 13317
rect 3973 13277 3985 13311
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 3050 13200 3056 13252
rect 3108 13240 3114 13252
rect 4080 13240 4108 13271
rect 4154 13268 4160 13320
rect 4212 13268 4218 13320
rect 5626 13268 5632 13320
rect 5684 13308 5690 13320
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 5684 13280 6009 13308
rect 5684 13268 5690 13280
rect 5997 13277 6009 13280
rect 6043 13308 6055 13311
rect 6546 13308 6552 13320
rect 6043 13280 6552 13308
rect 6043 13277 6055 13280
rect 5997 13271 6055 13277
rect 6546 13268 6552 13280
rect 6604 13268 6610 13320
rect 6638 13268 6644 13320
rect 6696 13268 6702 13320
rect 7116 13317 7144 13348
rect 7745 13345 7757 13348
rect 7791 13345 7803 13379
rect 7745 13339 7803 13345
rect 7966 13379 8024 13385
rect 7966 13345 7978 13379
rect 8012 13376 8024 13379
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 8012 13348 8493 13376
rect 8012 13345 8024 13348
rect 7966 13339 8024 13345
rect 8481 13345 8493 13348
rect 8527 13376 8539 13379
rect 9677 13379 9735 13385
rect 8527 13348 9536 13376
rect 8527 13345 8539 13348
rect 8481 13339 8539 13345
rect 9508 13320 9536 13348
rect 9677 13345 9689 13379
rect 9723 13376 9735 13379
rect 9950 13376 9956 13388
rect 9723 13348 9956 13376
rect 9723 13345 9735 13348
rect 9677 13339 9735 13345
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 7190 13268 7196 13320
rect 7248 13308 7254 13320
rect 7248 13280 8156 13308
rect 7248 13268 7254 13280
rect 8128 13252 8156 13280
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8567 13311 8625 13317
rect 8567 13308 8579 13311
rect 8260 13280 8579 13308
rect 8260 13268 8266 13280
rect 8567 13277 8579 13280
rect 8613 13308 8625 13311
rect 8613 13280 8800 13308
rect 8613 13277 8625 13280
rect 8567 13271 8625 13277
rect 5718 13240 5724 13252
rect 3108 13212 4108 13240
rect 4172 13212 5724 13240
rect 3108 13200 3114 13212
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 4172 13172 4200 13212
rect 5718 13200 5724 13212
rect 5776 13200 5782 13252
rect 7285 13243 7343 13249
rect 7285 13209 7297 13243
rect 7331 13240 7343 13243
rect 7331 13212 7788 13240
rect 7331 13209 7343 13212
rect 7285 13203 7343 13209
rect 3844 13144 4200 13172
rect 3844 13132 3850 13144
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 4304 13144 4353 13172
rect 4304 13132 4310 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 6270 13132 6276 13184
rect 6328 13132 6334 13184
rect 6914 13132 6920 13184
rect 6972 13132 6978 13184
rect 7466 13132 7472 13184
rect 7524 13132 7530 13184
rect 7760 13172 7788 13212
rect 8110 13200 8116 13252
rect 8168 13200 8174 13252
rect 8772 13240 8800 13280
rect 9490 13268 9496 13320
rect 9548 13308 9554 13320
rect 9585 13311 9643 13317
rect 9585 13308 9597 13311
rect 9548 13280 9597 13308
rect 9548 13268 9554 13280
rect 9585 13277 9597 13280
rect 9631 13277 9643 13311
rect 9585 13271 9643 13277
rect 10042 13240 10048 13252
rect 8772 13212 10048 13240
rect 10042 13200 10048 13212
rect 10100 13200 10106 13252
rect 7834 13172 7840 13184
rect 7760 13144 7840 13172
rect 7834 13132 7840 13144
rect 7892 13172 7898 13184
rect 8205 13175 8263 13181
rect 8205 13172 8217 13175
rect 7892 13144 8217 13172
rect 7892 13132 7898 13144
rect 8205 13141 8217 13144
rect 8251 13141 8263 13175
rect 8205 13135 8263 13141
rect 9674 13132 9680 13184
rect 9732 13172 9738 13184
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9732 13144 9965 13172
rect 9732 13132 9738 13144
rect 9953 13141 9965 13144
rect 9999 13172 10011 13175
rect 10410 13172 10416 13184
rect 9999 13144 10416 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 1104 13082 13340 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 13340 13082
rect 1104 13008 13340 13030
rect 4617 12971 4675 12977
rect 4617 12937 4629 12971
rect 4663 12968 4675 12971
rect 4982 12968 4988 12980
rect 4663 12940 4988 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 6914 12928 6920 12980
rect 6972 12928 6978 12980
rect 7190 12928 7196 12980
rect 7248 12928 7254 12980
rect 8297 12971 8355 12977
rect 8297 12968 8309 12971
rect 7392 12940 8309 12968
rect 6932 12900 6960 12928
rect 7392 12909 7420 12940
rect 8297 12937 8309 12940
rect 8343 12937 8355 12971
rect 9674 12968 9680 12980
rect 8297 12931 8355 12937
rect 8680 12940 9680 12968
rect 7377 12903 7435 12909
rect 3896 12872 4844 12900
rect 3786 12792 3792 12844
rect 3844 12792 3850 12844
rect 3896 12773 3924 12872
rect 4157 12835 4215 12841
rect 4157 12801 4169 12835
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12733 3939 12767
rect 4172 12764 4200 12795
rect 4246 12792 4252 12844
rect 4304 12792 4310 12844
rect 4433 12835 4491 12841
rect 4433 12801 4445 12835
rect 4479 12832 4491 12835
rect 4479 12804 4660 12832
rect 4479 12801 4491 12804
rect 4433 12795 4491 12801
rect 4522 12764 4528 12776
rect 4172 12736 4528 12764
rect 3881 12727 3939 12733
rect 4522 12724 4528 12736
rect 4580 12724 4586 12776
rect 4632 12764 4660 12804
rect 4706 12792 4712 12844
rect 4764 12792 4770 12844
rect 4632 12736 4752 12764
rect 4724 12708 4752 12736
rect 4338 12656 4344 12708
rect 4396 12656 4402 12708
rect 4706 12656 4712 12708
rect 4764 12656 4770 12708
rect 4816 12705 4844 12872
rect 6196 12872 6776 12900
rect 6932 12872 7328 12900
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 5258 12832 5264 12844
rect 5184 12804 5264 12832
rect 4985 12767 5043 12773
rect 4985 12733 4997 12767
rect 5031 12764 5043 12767
rect 5184 12764 5212 12804
rect 5258 12792 5264 12804
rect 5316 12792 5322 12844
rect 5537 12835 5595 12841
rect 5537 12801 5549 12835
rect 5583 12832 5595 12835
rect 5626 12832 5632 12844
rect 5583 12804 5632 12832
rect 5583 12801 5595 12804
rect 5537 12795 5595 12801
rect 5626 12792 5632 12804
rect 5684 12792 5690 12844
rect 6196 12841 6224 12872
rect 6181 12835 6239 12841
rect 6181 12801 6193 12835
rect 6227 12801 6239 12835
rect 6181 12795 6239 12801
rect 6546 12792 6552 12844
rect 6604 12832 6610 12844
rect 6641 12835 6699 12841
rect 6641 12832 6653 12835
rect 6604 12804 6653 12832
rect 6604 12792 6610 12804
rect 6641 12801 6653 12804
rect 6687 12801 6699 12835
rect 6748 12832 6776 12872
rect 6917 12835 6975 12841
rect 6917 12832 6929 12835
rect 6748 12804 6929 12832
rect 6641 12795 6699 12801
rect 6917 12801 6929 12804
rect 6963 12801 6975 12835
rect 6917 12795 6975 12801
rect 5031 12736 5212 12764
rect 5399 12767 5457 12773
rect 5031 12733 5043 12736
rect 4985 12727 5043 12733
rect 5399 12733 5411 12767
rect 5445 12764 5457 12767
rect 6822 12764 6828 12776
rect 5445 12736 6828 12764
rect 5445 12733 5457 12736
rect 5399 12727 5457 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 6932 12764 6960 12795
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7300 12841 7328 12872
rect 7377 12869 7389 12903
rect 7423 12869 7435 12903
rect 7377 12863 7435 12869
rect 7561 12903 7619 12909
rect 7561 12869 7573 12903
rect 7607 12900 7619 12903
rect 8481 12903 8539 12909
rect 8481 12900 8493 12903
rect 7607 12872 8493 12900
rect 7607 12869 7619 12872
rect 7561 12863 7619 12869
rect 8481 12869 8493 12872
rect 8527 12869 8539 12903
rect 8481 12863 8539 12869
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 7650 12792 7656 12844
rect 7708 12792 7714 12844
rect 7742 12792 7748 12844
rect 7800 12792 7806 12844
rect 8680 12841 8708 12940
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 9950 12928 9956 12980
rect 10008 12968 10014 12980
rect 10008 12940 10180 12968
rect 10008 12928 10014 12940
rect 9490 12900 9496 12912
rect 9140 12872 9496 12900
rect 7929 12835 7987 12841
rect 7929 12801 7941 12835
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12801 8079 12835
rect 8021 12795 8079 12801
rect 8113 12835 8171 12841
rect 8113 12801 8125 12835
rect 8159 12801 8171 12835
rect 8113 12795 8171 12801
rect 8665 12835 8723 12841
rect 8665 12801 8677 12835
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12832 8815 12835
rect 8846 12832 8852 12844
rect 8803 12804 8852 12832
rect 8803 12801 8815 12804
rect 8757 12795 8815 12801
rect 7466 12764 7472 12776
rect 6932 12736 7472 12764
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 4801 12699 4859 12705
rect 4801 12665 4813 12699
rect 4847 12696 4859 12699
rect 6362 12696 6368 12708
rect 4847 12668 6368 12696
rect 4847 12665 4859 12668
rect 4801 12659 4859 12665
rect 6362 12656 6368 12668
rect 6420 12696 6426 12708
rect 6457 12699 6515 12705
rect 6457 12696 6469 12699
rect 6420 12668 6469 12696
rect 6420 12656 6426 12668
rect 6457 12665 6469 12668
rect 6503 12665 6515 12699
rect 6457 12659 6515 12665
rect 7374 12656 7380 12708
rect 7432 12656 7438 12708
rect 3510 12588 3516 12640
rect 3568 12588 3574 12640
rect 4893 12631 4951 12637
rect 4893 12597 4905 12631
rect 4939 12628 4951 12631
rect 5074 12628 5080 12640
rect 4939 12600 5080 12628
rect 4939 12597 4951 12600
rect 4893 12591 4951 12597
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 5166 12588 5172 12640
rect 5224 12588 5230 12640
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5721 12631 5779 12637
rect 5721 12628 5733 12631
rect 5307 12600 5733 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5721 12597 5733 12600
rect 5767 12597 5779 12631
rect 5721 12591 5779 12597
rect 6730 12588 6736 12640
rect 6788 12588 6794 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7009 12631 7067 12637
rect 7009 12628 7021 12631
rect 6972 12600 7021 12628
rect 6972 12588 6978 12600
rect 7009 12597 7021 12600
rect 7055 12628 7067 12631
rect 7944 12628 7972 12795
rect 8036 12696 8064 12795
rect 8128 12764 8156 12795
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9140 12841 9168 12872
rect 9490 12860 9496 12872
rect 9548 12860 9554 12912
rect 10152 12909 10180 12940
rect 10137 12903 10195 12909
rect 10137 12869 10149 12903
rect 10183 12869 10195 12903
rect 10137 12863 10195 12869
rect 10612 12872 10916 12900
rect 9033 12835 9091 12841
rect 9033 12801 9045 12835
rect 9079 12801 9091 12835
rect 9033 12795 9091 12801
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12801 9183 12835
rect 9125 12795 9183 12801
rect 8294 12764 8300 12776
rect 8128 12736 8300 12764
rect 8294 12724 8300 12736
rect 8352 12764 8358 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8352 12736 8953 12764
rect 8352 12724 8358 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 8386 12696 8392 12708
rect 8036 12668 8392 12696
rect 8386 12656 8392 12668
rect 8444 12696 8450 12708
rect 9048 12696 9076 12795
rect 9398 12792 9404 12844
rect 9456 12792 9462 12844
rect 9858 12792 9864 12844
rect 9916 12792 9922 12844
rect 10042 12792 10048 12844
rect 10100 12832 10106 12844
rect 10612 12832 10640 12872
rect 10888 12841 10916 12872
rect 10100 12804 10640 12832
rect 10689 12835 10747 12841
rect 10100 12792 10106 12804
rect 10689 12801 10701 12835
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 11238 12832 11244 12844
rect 10919 12804 11244 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 9876 12764 9904 12792
rect 10704 12764 10732 12795
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 9876 12736 10732 12764
rect 8444 12668 9076 12696
rect 10505 12699 10563 12705
rect 8444 12656 8450 12668
rect 10505 12665 10517 12699
rect 10551 12696 10563 12699
rect 10781 12699 10839 12705
rect 10781 12696 10793 12699
rect 10551 12668 10793 12696
rect 10551 12665 10563 12668
rect 10505 12659 10563 12665
rect 10781 12665 10793 12668
rect 10827 12665 10839 12699
rect 10781 12659 10839 12665
rect 7055 12600 7972 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 9214 12588 9220 12640
rect 9272 12588 9278 12640
rect 9490 12588 9496 12640
rect 9548 12588 9554 12640
rect 10594 12588 10600 12640
rect 10652 12588 10658 12640
rect 1104 12538 13340 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 13340 12538
rect 1104 12464 13340 12486
rect 3050 12384 3056 12436
rect 3108 12384 3114 12436
rect 3513 12427 3571 12433
rect 3513 12393 3525 12427
rect 3559 12424 3571 12427
rect 3602 12424 3608 12436
rect 3559 12396 3608 12424
rect 3559 12393 3571 12396
rect 3513 12387 3571 12393
rect 3602 12384 3608 12396
rect 3660 12384 3666 12436
rect 4062 12384 4068 12436
rect 4120 12384 4126 12436
rect 5905 12427 5963 12433
rect 5905 12393 5917 12427
rect 5951 12424 5963 12427
rect 6270 12424 6276 12436
rect 5951 12396 6276 12424
rect 5951 12393 5963 12396
rect 5905 12387 5963 12393
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 6917 12427 6975 12433
rect 6917 12393 6929 12427
rect 6963 12424 6975 12427
rect 7006 12424 7012 12436
rect 6963 12396 7012 12424
rect 6963 12393 6975 12396
rect 6917 12387 6975 12393
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 11330 12384 11336 12436
rect 11388 12384 11394 12436
rect 6016 12359 6074 12365
rect 6016 12325 6028 12359
rect 6062 12356 6074 12359
rect 6062 12328 6132 12356
rect 6062 12325 6074 12328
rect 6016 12319 6074 12325
rect 3786 12288 3792 12300
rect 3344 12260 3792 12288
rect 3344 12229 3372 12260
rect 3786 12248 3792 12260
rect 3844 12248 3850 12300
rect 4338 12288 4344 12300
rect 4172 12260 4344 12288
rect 3237 12223 3295 12229
rect 3237 12189 3249 12223
rect 3283 12189 3295 12223
rect 3237 12183 3295 12189
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3605 12223 3663 12229
rect 3605 12189 3617 12223
rect 3651 12220 3663 12223
rect 4172 12220 4200 12260
rect 4338 12248 4344 12260
rect 4396 12248 4402 12300
rect 4522 12248 4528 12300
rect 4580 12248 4586 12300
rect 5074 12288 5080 12300
rect 4632 12260 5080 12288
rect 3651 12192 4200 12220
rect 3651 12189 3663 12192
rect 3605 12183 3663 12189
rect 3252 12152 3280 12183
rect 4246 12180 4252 12232
rect 4304 12180 4310 12232
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4632 12231 4660 12260
rect 5074 12248 5080 12260
rect 5132 12248 5138 12300
rect 5813 12291 5871 12297
rect 5813 12257 5825 12291
rect 5859 12288 5871 12291
rect 5902 12288 5908 12300
rect 5859 12260 5908 12288
rect 5859 12257 5871 12260
rect 5813 12251 5871 12257
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 4617 12225 4675 12231
rect 4617 12191 4629 12225
rect 4663 12191 4675 12225
rect 4801 12223 4859 12229
rect 4801 12198 4813 12223
rect 4617 12185 4675 12191
rect 4724 12189 4813 12198
rect 4847 12189 4859 12223
rect 4724 12183 4859 12189
rect 4724 12170 4844 12183
rect 3510 12152 3516 12164
rect 3252 12124 3516 12152
rect 3510 12112 3516 12124
rect 3568 12112 3574 12164
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4724 12152 4752 12170
rect 4212 12124 4752 12152
rect 6104 12152 6132 12328
rect 8294 12316 8300 12368
rect 8352 12316 8358 12368
rect 9122 12316 9128 12368
rect 9180 12356 9186 12368
rect 10597 12359 10655 12365
rect 9180 12328 9674 12356
rect 9180 12316 9186 12328
rect 7834 12248 7840 12300
rect 7892 12248 7898 12300
rect 8478 12288 8484 12300
rect 7944 12260 8484 12288
rect 6181 12223 6239 12229
rect 6181 12189 6193 12223
rect 6227 12220 6239 12223
rect 6733 12223 6791 12229
rect 6733 12220 6745 12223
rect 6227 12192 6745 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6733 12189 6745 12192
rect 6779 12220 6791 12223
rect 6822 12220 6828 12232
rect 6779 12192 6828 12220
rect 6779 12189 6791 12192
rect 6733 12183 6791 12189
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 6917 12223 6975 12229
rect 6917 12189 6929 12223
rect 6963 12220 6975 12223
rect 7466 12220 7472 12232
rect 6963 12192 7472 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 6932 12152 6960 12183
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7944 12229 7972 12260
rect 8478 12248 8484 12260
rect 8536 12288 8542 12300
rect 9646 12288 9674 12328
rect 10597 12325 10609 12359
rect 10643 12356 10655 12359
rect 10643 12328 11284 12356
rect 10643 12325 10655 12328
rect 10597 12319 10655 12325
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 8536 12260 9536 12288
rect 9646 12260 10088 12288
rect 8536 12248 8542 12260
rect 9508 12232 9536 12260
rect 10060 12232 10088 12260
rect 10244 12260 10793 12288
rect 7929 12223 7987 12229
rect 7929 12189 7941 12223
rect 7975 12189 7987 12223
rect 7929 12183 7987 12189
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 8168 12192 8401 12220
rect 8168 12180 8174 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 8570 12180 8576 12232
rect 8628 12220 8634 12232
rect 9122 12220 9128 12232
rect 8628 12192 9128 12220
rect 8628 12180 8634 12192
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 9490 12180 9496 12232
rect 9548 12180 9554 12232
rect 9769 12223 9827 12229
rect 9769 12189 9781 12223
rect 9815 12220 9827 12223
rect 9858 12220 9864 12232
rect 9815 12192 9864 12220
rect 9815 12189 9827 12192
rect 9769 12183 9827 12189
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 10244 12229 10272 12260
rect 10612 12232 10640 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 10229 12223 10287 12229
rect 10229 12189 10241 12223
rect 10275 12189 10287 12223
rect 10229 12183 10287 12189
rect 10410 12180 10416 12232
rect 10468 12180 10474 12232
rect 10594 12180 10600 12232
rect 10652 12180 10658 12232
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 6104 12124 6960 12152
rect 9309 12155 9367 12161
rect 4212 12112 4218 12124
rect 9309 12121 9321 12155
rect 9355 12152 9367 12155
rect 9950 12152 9956 12164
rect 9355 12124 9956 12152
rect 9355 12121 9367 12124
rect 9309 12115 9367 12121
rect 3326 12044 3332 12096
rect 3384 12084 3390 12096
rect 4430 12084 4436 12096
rect 3384 12056 4436 12084
rect 3384 12044 3390 12056
rect 4430 12044 4436 12056
rect 4488 12084 4494 12096
rect 5350 12084 5356 12096
rect 4488 12056 5356 12084
rect 4488 12044 4494 12056
rect 5350 12044 5356 12056
rect 5408 12044 5414 12096
rect 5537 12087 5595 12093
rect 5537 12053 5549 12087
rect 5583 12084 5595 12087
rect 5902 12084 5908 12096
rect 5583 12056 5908 12084
rect 5583 12053 5595 12056
rect 5537 12047 5595 12053
rect 5902 12044 5908 12056
rect 5960 12044 5966 12096
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 8481 12087 8539 12093
rect 8481 12084 8493 12087
rect 7984 12056 8493 12084
rect 7984 12044 7990 12056
rect 8481 12053 8493 12056
rect 8527 12053 8539 12087
rect 8481 12047 8539 12053
rect 8941 12087 8999 12093
rect 8941 12053 8953 12087
rect 8987 12084 8999 12087
rect 9030 12084 9036 12096
rect 8987 12056 9036 12084
rect 8987 12053 8999 12056
rect 8941 12047 8999 12053
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9122 12044 9128 12096
rect 9180 12084 9186 12096
rect 9324 12084 9352 12115
rect 9950 12112 9956 12124
rect 10008 12112 10014 12164
rect 10134 12112 10140 12164
rect 10192 12152 10198 12164
rect 10321 12155 10379 12161
rect 10321 12152 10333 12155
rect 10192 12124 10333 12152
rect 10192 12112 10198 12124
rect 10321 12121 10333 12124
rect 10367 12121 10379 12155
rect 10321 12115 10379 12121
rect 9180 12056 9352 12084
rect 9180 12044 9186 12056
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 9548 12056 9689 12084
rect 9548 12044 9554 12056
rect 9677 12053 9689 12056
rect 9723 12053 9735 12087
rect 9677 12047 9735 12053
rect 10042 12044 10048 12096
rect 10100 12084 10106 12096
rect 10704 12084 10732 12183
rect 10870 12180 10876 12232
rect 10928 12220 10934 12232
rect 10965 12223 11023 12229
rect 10965 12220 10977 12223
rect 10928 12192 10977 12220
rect 10928 12180 10934 12192
rect 10965 12189 10977 12192
rect 11011 12189 11023 12223
rect 10965 12183 11023 12189
rect 11054 12180 11060 12232
rect 11112 12180 11118 12232
rect 11256 12220 11284 12328
rect 11517 12223 11575 12229
rect 11517 12220 11529 12223
rect 11256 12192 11529 12220
rect 11517 12189 11529 12192
rect 11563 12189 11575 12223
rect 11517 12183 11575 12189
rect 11790 12180 11796 12232
rect 11848 12180 11854 12232
rect 10100 12056 10732 12084
rect 11241 12087 11299 12093
rect 10100 12044 10106 12056
rect 11241 12053 11253 12087
rect 11287 12084 11299 12087
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11287 12056 11713 12084
rect 11287 12053 11299 12056
rect 11241 12047 11299 12053
rect 11701 12053 11713 12056
rect 11747 12053 11759 12087
rect 11701 12047 11759 12053
rect 1104 11994 13340 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 13340 11994
rect 1104 11920 13340 11942
rect 4246 11880 4252 11892
rect 3252 11852 4252 11880
rect 3252 11753 3280 11852
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 4890 11880 4896 11892
rect 4396 11852 4896 11880
rect 4396 11840 4402 11852
rect 4890 11840 4896 11852
rect 4948 11880 4954 11892
rect 4948 11852 5120 11880
rect 4948 11840 4954 11852
rect 3510 11772 3516 11824
rect 3568 11812 3574 11824
rect 4264 11812 4292 11840
rect 4982 11812 4988 11824
rect 3568 11784 4108 11812
rect 4264 11784 4988 11812
rect 3568 11772 3574 11784
rect 4080 11756 4108 11784
rect 4982 11772 4988 11784
rect 5040 11772 5046 11824
rect 5092 11812 5120 11852
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5776 11852 6469 11880
rect 5776 11840 5782 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11790 11880 11796 11892
rect 11563 11852 11796 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12329 11883 12387 11889
rect 12329 11849 12341 11883
rect 12375 11880 12387 11883
rect 12618 11880 12624 11892
rect 12375 11852 12624 11880
rect 12375 11849 12387 11852
rect 12329 11843 12387 11849
rect 12618 11840 12624 11852
rect 12676 11840 12682 11892
rect 5092 11784 5396 11812
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11713 3295 11747
rect 3237 11707 3295 11713
rect 3786 11704 3792 11756
rect 3844 11744 3850 11756
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3844 11716 3985 11744
rect 3844 11704 3850 11716
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4062 11704 4068 11756
rect 4120 11704 4126 11756
rect 4154 11704 4160 11756
rect 4212 11704 4218 11756
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4798 11744 4804 11756
rect 4387 11716 4804 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4798 11704 4804 11716
rect 4856 11744 4862 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4856 11716 4905 11744
rect 4856 11704 4862 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5074 11704 5080 11756
rect 5132 11704 5138 11756
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11713 5227 11747
rect 5169 11707 5227 11713
rect 3326 11636 3332 11688
rect 3384 11636 3390 11688
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3697 11679 3755 11685
rect 3697 11676 3709 11679
rect 3467 11648 3709 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3697 11645 3709 11648
rect 3743 11645 3755 11679
rect 3697 11639 3755 11645
rect 5184 11620 5212 11707
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 5368 11753 5396 11784
rect 5902 11772 5908 11824
rect 5960 11772 5966 11824
rect 8478 11812 8484 11824
rect 8220 11784 8484 11812
rect 5368 11747 5437 11753
rect 5368 11716 5391 11747
rect 5379 11713 5391 11716
rect 5425 11713 5437 11747
rect 5379 11707 5437 11713
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 5684 11716 5825 11744
rect 5684 11704 5690 11716
rect 5813 11713 5825 11716
rect 5859 11713 5871 11747
rect 5920 11744 5948 11772
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5920 11716 6009 11744
rect 5813 11707 5871 11713
rect 5997 11713 6009 11716
rect 6043 11744 6055 11747
rect 6178 11744 6184 11756
rect 6043 11716 6184 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 6178 11704 6184 11716
rect 6236 11704 6242 11756
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11744 6423 11747
rect 6638 11744 6644 11756
rect 6411 11716 6644 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 7926 11704 7932 11756
rect 7984 11704 7990 11756
rect 8220 11753 8248 11784
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 12526 11772 12532 11824
rect 12584 11772 12590 11824
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11744 8355 11747
rect 8846 11744 8852 11756
rect 8343 11716 8852 11744
rect 8343 11713 8355 11716
rect 8297 11707 8355 11713
rect 8846 11704 8852 11716
rect 8904 11744 8910 11756
rect 9122 11744 9128 11756
rect 8904 11716 9128 11744
rect 8904 11704 8910 11716
rect 9122 11704 9128 11716
rect 9180 11704 9186 11756
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 5537 11679 5595 11685
rect 5537 11645 5549 11679
rect 5583 11676 5595 11679
rect 6454 11676 6460 11688
rect 5583 11648 6460 11676
rect 5583 11645 5595 11648
rect 5537 11639 5595 11645
rect 6454 11636 6460 11648
rect 6512 11636 6518 11688
rect 8021 11679 8079 11685
rect 8021 11645 8033 11679
rect 8067 11676 8079 11679
rect 8386 11676 8392 11688
rect 8067 11648 8392 11676
rect 8067 11645 8079 11648
rect 8021 11639 8079 11645
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 8570 11636 8576 11688
rect 8628 11676 8634 11688
rect 9232 11676 9260 11707
rect 9306 11704 9312 11756
rect 9364 11704 9370 11756
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11744 9643 11747
rect 9674 11744 9680 11756
rect 9631 11716 9680 11744
rect 9631 11713 9643 11716
rect 9585 11707 9643 11713
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11112 11716 11713 11744
rect 11112 11704 11118 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11793 11707 11851 11713
rect 8628 11648 9260 11676
rect 8628 11636 8634 11648
rect 9490 11636 9496 11688
rect 9548 11636 9554 11688
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 11808 11676 11836 11707
rect 11882 11704 11888 11756
rect 11940 11704 11946 11756
rect 12066 11704 12072 11756
rect 12124 11704 12130 11756
rect 10928 11648 11836 11676
rect 10928 11636 10934 11648
rect 3605 11611 3663 11617
rect 3605 11577 3617 11611
rect 3651 11608 3663 11611
rect 4706 11608 4712 11620
rect 3651 11580 4712 11608
rect 3651 11577 3663 11580
rect 3605 11571 3663 11577
rect 4706 11568 4712 11580
rect 4764 11568 4770 11620
rect 5166 11568 5172 11620
rect 5224 11608 5230 11620
rect 6362 11608 6368 11620
rect 5224 11580 6368 11608
rect 5224 11568 5230 11580
rect 6362 11568 6368 11580
rect 6420 11568 6426 11620
rect 3421 11543 3479 11549
rect 3421 11509 3433 11543
rect 3467 11540 3479 11543
rect 4614 11540 4620 11552
rect 3467 11512 4620 11540
rect 3467 11509 3479 11512
rect 3421 11503 3479 11509
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 5350 11500 5356 11552
rect 5408 11540 5414 11552
rect 5626 11540 5632 11552
rect 5408 11512 5632 11540
rect 5408 11500 5414 11512
rect 5626 11500 5632 11512
rect 5684 11500 5690 11552
rect 8478 11500 8484 11552
rect 8536 11500 8542 11552
rect 8938 11500 8944 11552
rect 8996 11540 9002 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8996 11512 9045 11540
rect 8996 11500 9002 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 9033 11503 9091 11509
rect 12161 11543 12219 11549
rect 12161 11509 12173 11543
rect 12207 11540 12219 11543
rect 12250 11540 12256 11552
rect 12207 11512 12256 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12345 11543 12403 11549
rect 12345 11509 12357 11543
rect 12391 11540 12403 11543
rect 12710 11540 12716 11552
rect 12391 11512 12716 11540
rect 12391 11509 12403 11512
rect 12345 11503 12403 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 1104 11450 13340 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 13340 11450
rect 1104 11376 13340 11398
rect 3881 11339 3939 11345
rect 3881 11305 3893 11339
rect 3927 11336 3939 11339
rect 4062 11336 4068 11348
rect 3927 11308 4068 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4433 11339 4491 11345
rect 4433 11305 4445 11339
rect 4479 11336 4491 11339
rect 4706 11336 4712 11348
rect 4479 11308 4712 11336
rect 4479 11305 4491 11308
rect 4433 11299 4491 11305
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 4948 11308 5856 11336
rect 4948 11296 4954 11308
rect 5166 11268 5172 11280
rect 4264 11240 5172 11268
rect 4264 11141 4292 11240
rect 5166 11228 5172 11240
rect 5224 11228 5230 11280
rect 5074 11200 5080 11212
rect 4356 11172 5080 11200
rect 4356 11141 4384 11172
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 5626 11200 5632 11212
rect 5184 11172 5632 11200
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3896 11104 4077 11132
rect 3510 10956 3516 11008
rect 3568 10996 3574 11008
rect 3896 10996 3924 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 4632 11064 4660 11095
rect 4982 11092 4988 11144
rect 5040 11092 5046 11144
rect 5184 11132 5212 11172
rect 5626 11160 5632 11172
rect 5684 11160 5690 11212
rect 5828 11141 5856 11308
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11517 11339 11575 11345
rect 11517 11336 11529 11339
rect 11112 11308 11529 11336
rect 11112 11296 11118 11308
rect 11517 11305 11529 11308
rect 11563 11305 11575 11339
rect 11517 11299 11575 11305
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8481 11203 8539 11209
rect 8481 11200 8493 11203
rect 7984 11172 8493 11200
rect 7984 11160 7990 11172
rect 8481 11169 8493 11172
rect 8527 11169 8539 11203
rect 8481 11163 8539 11169
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11333 11203 11391 11209
rect 11333 11200 11345 11203
rect 11296 11172 11345 11200
rect 11296 11160 11302 11172
rect 11333 11169 11345 11172
rect 11379 11169 11391 11203
rect 12710 11200 12716 11212
rect 11333 11163 11391 11169
rect 11808 11172 12716 11200
rect 5092 11104 5212 11132
rect 5537 11135 5595 11141
rect 4028 11036 4660 11064
rect 4028 11024 4034 11036
rect 4706 11024 4712 11076
rect 4764 11024 4770 11076
rect 4801 11067 4859 11073
rect 4801 11033 4813 11067
rect 4847 11064 4859 11067
rect 5092 11064 5120 11104
rect 5537 11101 5549 11135
rect 5583 11101 5595 11135
rect 5537 11095 5595 11101
rect 5813 11135 5871 11141
rect 5813 11101 5825 11135
rect 5859 11101 5871 11135
rect 5813 11095 5871 11101
rect 8297 11135 8355 11141
rect 8297 11101 8309 11135
rect 8343 11132 8355 11135
rect 8386 11132 8392 11144
rect 8343 11104 8392 11132
rect 8343 11101 8355 11104
rect 8297 11095 8355 11101
rect 4847 11036 5120 11064
rect 5552 11064 5580 11095
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11132 9459 11135
rect 9490 11132 9496 11144
rect 9447 11104 9496 11132
rect 9447 11101 9459 11104
rect 9401 11095 9459 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 9674 11132 9680 11144
rect 9631 11104 9680 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 9674 11092 9680 11104
rect 9732 11132 9738 11144
rect 10870 11132 10876 11144
rect 9732 11104 10876 11132
rect 9732 11092 9738 11104
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 11808 11141 11836 11172
rect 12710 11160 12716 11172
rect 12768 11160 12774 11212
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12802 11132 12808 11144
rect 12207 11104 12808 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12802 11092 12808 11104
rect 12860 11092 12866 11144
rect 12894 11092 12900 11144
rect 12952 11092 12958 11144
rect 6270 11064 6276 11076
rect 5552 11036 6276 11064
rect 4847 11033 4859 11036
rect 4801 11027 4859 11033
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 12434 11024 12440 11076
rect 12492 11024 12498 11076
rect 5258 10996 5264 11008
rect 3568 10968 5264 10996
rect 3568 10956 3574 10968
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 5442 10956 5448 11008
rect 5500 10956 5506 11008
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8113 10999 8171 11005
rect 8113 10996 8125 10999
rect 8076 10968 8125 10996
rect 8076 10956 8082 10968
rect 8113 10965 8125 10968
rect 8159 10965 8171 10999
rect 8113 10959 8171 10965
rect 9490 10956 9496 11008
rect 9548 10956 9554 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 11701 10999 11759 11005
rect 11701 10996 11713 10999
rect 10376 10968 11713 10996
rect 10376 10956 10382 10968
rect 11701 10965 11713 10968
rect 11747 10996 11759 10999
rect 11974 10996 11980 11008
rect 11747 10968 11980 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 1104 10906 13340 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 13340 10906
rect 1104 10832 13340 10854
rect 11882 10752 11888 10804
rect 11940 10792 11946 10804
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 11940 10764 12357 10792
rect 11940 10752 11946 10764
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12345 10755 12403 10761
rect 3878 10724 3884 10736
rect 2806 10696 3884 10724
rect 3878 10684 3884 10696
rect 3936 10684 3942 10736
rect 5902 10684 5908 10736
rect 5960 10724 5966 10736
rect 5997 10727 6055 10733
rect 5997 10724 6009 10727
rect 5960 10696 6009 10724
rect 5960 10684 5966 10696
rect 5997 10693 6009 10696
rect 6043 10693 6055 10727
rect 5997 10687 6055 10693
rect 8205 10727 8263 10733
rect 8205 10693 8217 10727
rect 8251 10724 8263 10727
rect 8478 10724 8484 10736
rect 8251 10696 8484 10724
rect 8251 10693 8263 10696
rect 8205 10687 8263 10693
rect 5258 10616 5264 10668
rect 5316 10656 5322 10668
rect 5534 10656 5540 10668
rect 5316 10628 5540 10656
rect 5316 10616 5322 10628
rect 5534 10616 5540 10628
rect 5592 10616 5598 10668
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10656 5687 10659
rect 5718 10656 5724 10668
rect 5675 10628 5724 10656
rect 5675 10625 5687 10628
rect 5629 10619 5687 10625
rect 5718 10616 5724 10628
rect 5776 10616 5782 10668
rect 1489 10591 1547 10597
rect 1489 10557 1501 10591
rect 1535 10588 1547 10591
rect 1670 10588 1676 10600
rect 1535 10560 1676 10588
rect 1535 10557 1547 10560
rect 1489 10551 1547 10557
rect 1670 10548 1676 10560
rect 1728 10548 1734 10600
rect 3234 10548 3240 10600
rect 3292 10548 3298 10600
rect 3513 10591 3571 10597
rect 3513 10557 3525 10591
rect 3559 10557 3571 10591
rect 3513 10551 3571 10557
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3528 10452 3556 10551
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 5905 10591 5963 10597
rect 5905 10588 5917 10591
rect 5868 10560 5917 10588
rect 5868 10548 5874 10560
rect 5905 10557 5917 10560
rect 5951 10557 5963 10591
rect 6012 10588 6040 10687
rect 8478 10684 8484 10696
rect 8536 10724 8542 10736
rect 9214 10724 9220 10736
rect 8536 10696 9220 10724
rect 8536 10684 8542 10696
rect 9214 10684 9220 10696
rect 9272 10684 9278 10736
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 11517 10727 11575 10733
rect 11517 10724 11529 10727
rect 11296 10696 11529 10724
rect 11296 10684 11302 10696
rect 11517 10693 11529 10696
rect 11563 10693 11575 10727
rect 11517 10687 11575 10693
rect 11974 10684 11980 10736
rect 12032 10724 12038 10736
rect 12253 10727 12311 10733
rect 12253 10724 12265 10727
rect 12032 10696 12265 10724
rect 12032 10684 12038 10696
rect 12253 10693 12265 10696
rect 12299 10693 12311 10727
rect 12253 10687 12311 10693
rect 12618 10684 12624 10736
rect 12676 10724 12682 10736
rect 12676 10696 12848 10724
rect 12676 10684 12682 10696
rect 12820 10668 12848 10696
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6917 10659 6975 10665
rect 6604 10628 6868 10656
rect 6604 10616 6610 10628
rect 6840 10597 6868 10628
rect 6917 10625 6929 10659
rect 6963 10656 6975 10659
rect 7466 10656 7472 10668
rect 6963 10628 7472 10656
rect 6963 10625 6975 10628
rect 6917 10619 6975 10625
rect 7466 10616 7472 10628
rect 7524 10616 7530 10668
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 8297 10619 8355 10625
rect 6733 10591 6791 10597
rect 6733 10588 6745 10591
rect 6012 10560 6745 10588
rect 5905 10551 5963 10557
rect 6733 10557 6745 10560
rect 6779 10557 6791 10591
rect 6733 10551 6791 10557
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10588 6883 10591
rect 7374 10588 7380 10600
rect 6871 10560 7380 10588
rect 6871 10557 6883 10560
rect 6825 10551 6883 10557
rect 5920 10520 5948 10551
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 8312 10588 8340 10619
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9030 10616 9036 10668
rect 9088 10616 9094 10668
rect 9306 10616 9312 10668
rect 9364 10656 9370 10668
rect 9490 10656 9496 10668
rect 9364 10628 9496 10656
rect 9364 10616 9370 10628
rect 9490 10616 9496 10628
rect 9548 10616 9554 10668
rect 9674 10616 9680 10668
rect 9732 10616 9738 10668
rect 12526 10656 12532 10668
rect 10980 10628 12532 10656
rect 8573 10591 8631 10597
rect 8573 10588 8585 10591
rect 8312 10560 8585 10588
rect 8573 10557 8585 10560
rect 8619 10557 8631 10591
rect 8573 10551 8631 10557
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 6549 10523 6607 10529
rect 6549 10520 6561 10523
rect 5920 10492 6561 10520
rect 6549 10489 6561 10492
rect 6595 10489 6607 10523
rect 8772 10520 8800 10551
rect 8846 10548 8852 10600
rect 8904 10548 8910 10600
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 10318 10548 10324 10600
rect 10376 10548 10382 10600
rect 9217 10523 9275 10529
rect 9217 10520 9229 10523
rect 8772 10492 9229 10520
rect 6549 10483 6607 10489
rect 9217 10489 9229 10492
rect 9263 10489 9275 10523
rect 9217 10483 9275 10489
rect 10045 10523 10103 10529
rect 10045 10489 10057 10523
rect 10091 10520 10103 10523
rect 10226 10520 10232 10532
rect 10091 10492 10232 10520
rect 10091 10489 10103 10492
rect 10045 10483 10103 10489
rect 10226 10480 10232 10492
rect 10284 10520 10290 10532
rect 10980 10520 11008 10628
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 12710 10616 12716 10668
rect 12768 10616 12774 10668
rect 12802 10616 12808 10668
rect 12860 10616 12866 10668
rect 11885 10591 11943 10597
rect 11885 10557 11897 10591
rect 11931 10588 11943 10591
rect 12434 10588 12440 10600
rect 11931 10560 12440 10588
rect 11931 10557 11943 10560
rect 11885 10551 11943 10557
rect 12434 10548 12440 10560
rect 12492 10548 12498 10600
rect 10284 10492 11008 10520
rect 11977 10523 12035 10529
rect 10284 10480 10290 10492
rect 11977 10489 11989 10523
rect 12023 10520 12035 10523
rect 12526 10520 12532 10532
rect 12023 10492 12532 10520
rect 12023 10489 12035 10492
rect 11977 10483 12035 10489
rect 12526 10480 12532 10492
rect 12584 10480 12590 10532
rect 2832 10424 3556 10452
rect 5353 10455 5411 10461
rect 2832 10412 2838 10424
rect 5353 10421 5365 10455
rect 5399 10452 5411 10455
rect 6638 10452 6644 10464
rect 5399 10424 6644 10452
rect 5399 10421 5411 10424
rect 5353 10415 5411 10421
rect 6638 10412 6644 10424
rect 6696 10412 6702 10464
rect 6730 10412 6736 10464
rect 6788 10412 6794 10464
rect 7282 10412 7288 10464
rect 7340 10452 7346 10464
rect 7837 10455 7895 10461
rect 7837 10452 7849 10455
rect 7340 10424 7849 10452
rect 7340 10412 7346 10424
rect 7837 10421 7849 10424
rect 7883 10421 7895 10455
rect 7837 10415 7895 10421
rect 8110 10412 8116 10464
rect 8168 10452 8174 10464
rect 9582 10452 9588 10464
rect 8168 10424 9588 10452
rect 8168 10412 8174 10424
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9858 10412 9864 10464
rect 9916 10412 9922 10464
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 12115 10455 12173 10461
rect 12115 10452 12127 10455
rect 10744 10424 12127 10452
rect 10744 10412 10750 10424
rect 12115 10421 12127 10424
rect 12161 10452 12173 10455
rect 12618 10452 12624 10464
rect 12161 10424 12624 10452
rect 12161 10421 12173 10424
rect 12115 10415 12173 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 1104 10362 13340 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 13340 10362
rect 1104 10288 13340 10310
rect 3510 10208 3516 10260
rect 3568 10208 3574 10260
rect 3878 10208 3884 10260
rect 3936 10208 3942 10260
rect 4706 10208 4712 10260
rect 4764 10208 4770 10260
rect 6638 10208 6644 10260
rect 6696 10248 6702 10260
rect 9493 10251 9551 10257
rect 6696 10220 9352 10248
rect 6696 10208 6702 10220
rect 4724 10180 4752 10208
rect 7009 10183 7067 10189
rect 4264 10152 5396 10180
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 2774 10112 2780 10124
rect 1811 10084 2780 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3786 10112 3792 10124
rect 3108 10084 3792 10112
rect 3108 10072 3114 10084
rect 3786 10072 3792 10084
rect 3844 10112 3850 10124
rect 4264 10121 4292 10152
rect 5368 10121 5396 10152
rect 7009 10149 7021 10183
rect 7055 10149 7067 10183
rect 8665 10183 8723 10189
rect 8665 10180 8677 10183
rect 7009 10143 7067 10149
rect 7208 10152 8677 10180
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3844 10084 4261 10112
rect 3844 10072 3850 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 5353 10115 5411 10121
rect 4249 10075 4307 10081
rect 4356 10084 5304 10112
rect 1486 10004 1492 10056
rect 1544 10004 1550 10056
rect 1670 10004 1676 10056
rect 1728 10004 1734 10056
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10044 4031 10047
rect 4062 10044 4068 10056
rect 4019 10016 4068 10044
rect 4019 10013 4031 10016
rect 3973 10007 4031 10013
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4157 10047 4215 10053
rect 4157 10013 4169 10047
rect 4203 10044 4215 10047
rect 4356 10044 4384 10084
rect 4203 10016 4384 10044
rect 4433 10047 4491 10053
rect 4203 10013 4215 10016
rect 4157 10007 4215 10013
rect 4433 10013 4445 10047
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4706 10044 4712 10056
rect 4571 10016 4712 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 2038 9936 2044 9988
rect 2096 9936 2102 9988
rect 4448 9976 4476 10007
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 4798 10004 4804 10056
rect 4856 10004 4862 10056
rect 5276 10053 5304 10084
rect 5353 10081 5365 10115
rect 5399 10081 5411 10115
rect 7024 10112 7052 10143
rect 5353 10075 5411 10081
rect 6564 10084 7052 10112
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5442 10044 5448 10056
rect 5307 10016 5448 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 5442 10004 5448 10016
rect 5500 10004 5506 10056
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 5629 10047 5687 10053
rect 5629 10044 5641 10047
rect 5592 10016 5641 10044
rect 5592 10004 5598 10016
rect 5629 10013 5641 10016
rect 5675 10013 5687 10047
rect 5629 10007 5687 10013
rect 5718 10004 5724 10056
rect 5776 10004 5782 10056
rect 6564 10053 6592 10084
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10013 6331 10047
rect 6273 10007 6331 10013
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10013 6607 10047
rect 6549 10007 6607 10013
rect 4614 9976 4620 9988
rect 3266 9948 4200 9976
rect 4448 9948 4620 9976
rect 4172 9920 4200 9948
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 4985 9979 5043 9985
rect 4985 9945 4997 9979
rect 5031 9976 5043 9979
rect 5902 9976 5908 9988
rect 5031 9948 5908 9976
rect 5031 9945 5043 9948
rect 4985 9939 5043 9945
rect 5902 9936 5908 9948
rect 5960 9976 5966 9988
rect 6288 9976 6316 10007
rect 5960 9948 6316 9976
rect 5960 9936 5966 9948
rect 1673 9911 1731 9917
rect 1673 9877 1685 9911
rect 1719 9908 1731 9911
rect 3326 9908 3332 9920
rect 1719 9880 3332 9908
rect 1719 9877 1731 9880
rect 1673 9871 1731 9877
rect 3326 9868 3332 9880
rect 3384 9868 3390 9920
rect 4154 9868 4160 9920
rect 4212 9868 4218 9920
rect 4709 9911 4767 9917
rect 4709 9877 4721 9911
rect 4755 9908 4767 9911
rect 5534 9908 5540 9920
rect 4755 9880 5540 9908
rect 4755 9877 4767 9880
rect 4709 9871 4767 9877
rect 5534 9868 5540 9880
rect 5592 9908 5598 9920
rect 6472 9908 6500 10007
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 6730 10004 6736 10056
rect 6788 10044 6794 10056
rect 7009 10047 7067 10053
rect 7009 10044 7021 10047
rect 6788 10016 7021 10044
rect 6788 10004 6794 10016
rect 7009 10013 7021 10016
rect 7055 10044 7067 10047
rect 7208 10044 7236 10152
rect 8665 10149 8677 10152
rect 8711 10149 8723 10183
rect 8665 10143 8723 10149
rect 8754 10140 8760 10192
rect 8812 10180 8818 10192
rect 8941 10183 8999 10189
rect 8941 10180 8953 10183
rect 8812 10152 8953 10180
rect 8812 10140 8818 10152
rect 8941 10149 8953 10152
rect 8987 10149 8999 10183
rect 8941 10143 8999 10149
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 9217 10115 9275 10121
rect 9217 10112 9229 10115
rect 8076 10084 9229 10112
rect 8076 10072 8082 10084
rect 9217 10081 9229 10084
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 7055 10016 7236 10044
rect 7055 10013 7067 10016
rect 7009 10007 7067 10013
rect 7282 10004 7288 10056
rect 7340 10004 7346 10056
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7742 10044 7748 10056
rect 7515 10016 7748 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7742 10004 7748 10016
rect 7800 10004 7806 10056
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8938 10044 8944 10056
rect 8251 10016 8944 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 9324 10044 9352 10220
rect 9493 10217 9505 10251
rect 9539 10248 9551 10251
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 9539 10220 10333 10248
rect 9539 10217 9551 10220
rect 9493 10211 9551 10217
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 10321 10211 10379 10217
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 12434 10248 12440 10260
rect 10919 10220 12440 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 9582 10140 9588 10192
rect 9640 10180 9646 10192
rect 10413 10183 10471 10189
rect 10413 10180 10425 10183
rect 9640 10152 10425 10180
rect 9640 10140 9646 10152
rect 10413 10149 10425 10152
rect 10459 10149 10471 10183
rect 10413 10143 10471 10149
rect 10888 10112 10916 10211
rect 12434 10208 12440 10220
rect 12492 10208 12498 10260
rect 12710 10208 12716 10260
rect 12768 10248 12774 10260
rect 12805 10251 12863 10257
rect 12805 10248 12817 10251
rect 12768 10220 12817 10248
rect 12768 10208 12774 10220
rect 12805 10217 12817 10220
rect 12851 10217 12863 10251
rect 12805 10211 12863 10217
rect 11517 10183 11575 10189
rect 11517 10149 11529 10183
rect 11563 10149 11575 10183
rect 11517 10143 11575 10149
rect 11701 10183 11759 10189
rect 11701 10149 11713 10183
rect 11747 10180 11759 10183
rect 12066 10180 12072 10192
rect 11747 10152 12072 10180
rect 11747 10149 11759 10152
rect 11701 10143 11759 10149
rect 10520 10084 10916 10112
rect 9171 10016 9352 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 9674 10004 9680 10056
rect 9732 10004 9738 10056
rect 9766 10004 9772 10056
rect 9824 10004 9830 10056
rect 10183 10047 10241 10053
rect 10183 10013 10195 10047
rect 10229 10044 10241 10047
rect 10520 10044 10548 10084
rect 10229 10016 10548 10044
rect 10229 10013 10241 10016
rect 10183 10007 10241 10013
rect 10594 10004 10600 10056
rect 10652 10004 10658 10056
rect 10686 10004 10692 10056
rect 10744 10004 10750 10056
rect 10962 10044 10968 10056
rect 10796 10016 10968 10044
rect 7098 9936 7104 9988
rect 7156 9976 7162 9988
rect 7929 9979 7987 9985
rect 7929 9976 7941 9979
rect 7156 9948 7941 9976
rect 7156 9936 7162 9948
rect 7929 9945 7941 9948
rect 7975 9945 7987 9979
rect 7929 9939 7987 9945
rect 8665 9979 8723 9985
rect 8665 9945 8677 9979
rect 8711 9976 8723 9979
rect 9030 9976 9036 9988
rect 8711 9948 9036 9976
rect 8711 9945 8723 9948
rect 8665 9939 8723 9945
rect 9030 9936 9036 9948
rect 9088 9936 9094 9988
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 9585 9979 9643 9985
rect 9585 9976 9597 9979
rect 9272 9948 9597 9976
rect 9272 9936 9278 9948
rect 9585 9945 9597 9948
rect 9631 9945 9643 9979
rect 9585 9939 9643 9945
rect 9953 9979 10011 9985
rect 9953 9945 9965 9979
rect 9999 9945 10011 9979
rect 9953 9939 10011 9945
rect 10045 9979 10103 9985
rect 10045 9945 10057 9979
rect 10091 9976 10103 9979
rect 10796 9976 10824 10016
rect 10962 10004 10968 10016
rect 11020 10004 11026 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10044 11115 10047
rect 11238 10044 11244 10056
rect 11103 10016 11244 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11238 10004 11244 10016
rect 11296 10004 11302 10056
rect 11532 10044 11560 10143
rect 12066 10140 12072 10152
rect 12124 10140 12130 10192
rect 12526 10072 12532 10124
rect 12584 10072 12590 10124
rect 11839 10047 11897 10053
rect 11839 10044 11851 10047
rect 11532 10016 11851 10044
rect 11839 10013 11851 10016
rect 11885 10013 11897 10047
rect 11839 10007 11897 10013
rect 12158 10004 12164 10056
rect 12216 10053 12222 10056
rect 12216 10047 12255 10053
rect 12243 10013 12255 10047
rect 12216 10007 12255 10013
rect 12216 10004 12222 10007
rect 12342 10004 12348 10056
rect 12400 10004 12406 10056
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12618 10044 12624 10056
rect 12483 10016 12624 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 10091 9948 10824 9976
rect 10091 9945 10103 9948
rect 10045 9939 10103 9945
rect 5592 9880 6500 9908
rect 5592 9868 5598 9880
rect 6914 9868 6920 9920
rect 6972 9868 6978 9920
rect 7190 9868 7196 9920
rect 7248 9868 7254 9920
rect 7282 9868 7288 9920
rect 7340 9908 7346 9920
rect 7466 9908 7472 9920
rect 7340 9880 7472 9908
rect 7340 9868 7346 9880
rect 7466 9868 7472 9880
rect 7524 9908 7530 9920
rect 7561 9911 7619 9917
rect 7561 9908 7573 9911
rect 7524 9880 7573 9908
rect 7524 9868 7530 9880
rect 7561 9877 7573 9880
rect 7607 9908 7619 9911
rect 9968 9908 9996 9939
rect 11974 9936 11980 9988
rect 12032 9936 12038 9988
rect 12066 9936 12072 9988
rect 12124 9936 12130 9988
rect 7607 9880 9996 9908
rect 7607 9877 7619 9880
rect 7561 9871 7619 9877
rect 1104 9818 13340 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 13340 9818
rect 1104 9744 13340 9766
rect 2038 9664 2044 9716
rect 2096 9664 2102 9716
rect 2958 9704 2964 9716
rect 2148 9676 2964 9704
rect 1486 9596 1492 9648
rect 1544 9636 1550 9648
rect 1581 9639 1639 9645
rect 1581 9636 1593 9639
rect 1544 9608 1593 9636
rect 1544 9596 1550 9608
rect 1581 9605 1593 9608
rect 1627 9605 1639 9639
rect 1581 9599 1639 9605
rect 1596 9500 1624 9599
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 1765 9639 1823 9645
rect 1765 9636 1777 9639
rect 1728 9608 1777 9636
rect 1728 9596 1734 9608
rect 1765 9605 1777 9608
rect 1811 9636 1823 9639
rect 2148 9636 2176 9676
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 3234 9664 3240 9716
rect 3292 9704 3298 9716
rect 3605 9707 3663 9713
rect 3605 9704 3617 9707
rect 3292 9676 3617 9704
rect 3292 9664 3298 9676
rect 3605 9673 3617 9676
rect 3651 9673 3663 9707
rect 3605 9667 3663 9673
rect 4798 9664 4804 9716
rect 4856 9704 4862 9716
rect 4893 9707 4951 9713
rect 4893 9704 4905 9707
rect 4856 9676 4905 9704
rect 4856 9664 4862 9676
rect 4893 9673 4905 9676
rect 4939 9673 4951 9707
rect 7098 9704 7104 9716
rect 4893 9667 4951 9673
rect 6288 9676 7104 9704
rect 1811 9608 2176 9636
rect 2225 9639 2283 9645
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 2225 9605 2237 9639
rect 2271 9636 2283 9639
rect 2314 9636 2320 9648
rect 2271 9608 2320 9636
rect 2271 9605 2283 9608
rect 2225 9599 2283 9605
rect 2314 9596 2320 9608
rect 2372 9596 2378 9648
rect 3757 9639 3815 9645
rect 3757 9636 3769 9639
rect 2746 9608 3769 9636
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 2746 9568 2774 9608
rect 3757 9605 3769 9608
rect 3803 9605 3815 9639
rect 3757 9599 3815 9605
rect 3973 9639 4031 9645
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 4062 9636 4068 9648
rect 4019 9608 4068 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 4062 9596 4068 9608
rect 4120 9596 4126 9648
rect 4154 9596 4160 9648
rect 4212 9596 4218 9648
rect 1995 9540 2774 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 3108 9540 3341 9568
rect 3108 9528 3114 9540
rect 3329 9537 3341 9540
rect 3375 9568 3387 9571
rect 3878 9568 3884 9580
rect 3375 9540 3884 9568
rect 3375 9537 3387 9540
rect 3329 9531 3387 9537
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 4614 9528 4620 9580
rect 4672 9528 4678 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4798 9568 4804 9580
rect 4755 9540 4804 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 4908 9568 4936 9667
rect 5902 9596 5908 9648
rect 5960 9596 5966 9648
rect 6288 9636 6316 9676
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 7190 9664 7196 9716
rect 7248 9664 7254 9716
rect 8846 9664 8852 9716
rect 8904 9704 8910 9716
rect 9309 9707 9367 9713
rect 9309 9704 9321 9707
rect 8904 9676 9321 9704
rect 8904 9664 8910 9676
rect 9309 9673 9321 9676
rect 9355 9673 9367 9707
rect 9309 9667 9367 9673
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 10505 9707 10563 9713
rect 10505 9704 10517 9707
rect 9732 9676 10517 9704
rect 9732 9664 9738 9676
rect 10505 9673 10517 9676
rect 10551 9673 10563 9707
rect 10505 9667 10563 9673
rect 12066 9664 12072 9716
rect 12124 9664 12130 9716
rect 12526 9704 12532 9716
rect 12406 9676 12532 9704
rect 12406 9674 12434 9676
rect 6914 9636 6920 9648
rect 6012 9608 6316 9636
rect 6380 9608 6920 9636
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 4908 9540 5365 9568
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5534 9528 5540 9580
rect 5592 9568 5598 9580
rect 6012 9577 6040 9608
rect 5813 9571 5871 9577
rect 5813 9568 5825 9571
rect 5592 9540 5825 9568
rect 5592 9528 5598 9540
rect 5813 9537 5825 9540
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6086 9528 6092 9580
rect 6144 9528 6150 9580
rect 6380 9577 6408 9608
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 10226 9596 10232 9648
rect 10284 9596 10290 9648
rect 10594 9596 10600 9648
rect 10652 9636 10658 9648
rect 12268 9646 12434 9674
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 11149 9639 11207 9645
rect 11149 9636 11161 9639
rect 10652 9608 11161 9636
rect 10652 9596 10658 9608
rect 6365 9571 6423 9577
rect 6365 9537 6377 9571
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 6549 9571 6607 9577
rect 6549 9537 6561 9571
rect 6595 9568 6607 9571
rect 6595 9540 6776 9568
rect 6595 9537 6607 9540
rect 6549 9531 6607 9537
rect 2590 9500 2596 9512
rect 1596 9472 2596 9500
rect 2590 9460 2596 9472
rect 2648 9500 2654 9512
rect 3145 9503 3203 9509
rect 3145 9500 3157 9503
rect 2648 9472 3157 9500
rect 2648 9460 2654 9472
rect 3145 9469 3157 9472
rect 3191 9469 3203 9503
rect 3145 9463 3203 9469
rect 3510 9460 3516 9512
rect 3568 9460 3574 9512
rect 4264 9500 4292 9528
rect 5442 9500 5448 9512
rect 4264 9472 5448 9500
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9500 5687 9503
rect 6638 9500 6644 9512
rect 5675 9472 6644 9500
rect 5675 9469 5687 9472
rect 5629 9463 5687 9469
rect 6638 9460 6644 9472
rect 6696 9460 6702 9512
rect 2498 9392 2504 9444
rect 2556 9432 2562 9444
rect 2556 9404 2820 9432
rect 2556 9392 2562 9404
rect 2225 9367 2283 9373
rect 2225 9333 2237 9367
rect 2271 9364 2283 9367
rect 2685 9367 2743 9373
rect 2685 9364 2697 9367
rect 2271 9336 2697 9364
rect 2271 9333 2283 9336
rect 2225 9327 2283 9333
rect 2685 9333 2697 9336
rect 2731 9333 2743 9367
rect 2792 9364 2820 9404
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 3528 9432 3556 9460
rect 2924 9404 3556 9432
rect 5353 9435 5411 9441
rect 2924 9392 2930 9404
rect 5353 9401 5365 9435
rect 5399 9432 5411 9435
rect 6748 9432 6776 9540
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 7193 9571 7251 9577
rect 7193 9537 7205 9571
rect 7239 9568 7251 9571
rect 7282 9568 7288 9580
rect 7239 9540 7288 9568
rect 7239 9537 7251 9540
rect 7193 9531 7251 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7374 9528 7380 9580
rect 7432 9528 7438 9580
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9568 9275 9571
rect 9306 9568 9312 9580
rect 9263 9540 9312 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9568 9551 9571
rect 9539 9540 9812 9568
rect 9539 9537 9551 9540
rect 9493 9531 9551 9537
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9508 9500 9536 9531
rect 9784 9509 9812 9540
rect 10686 9528 10692 9580
rect 10744 9528 10750 9580
rect 10796 9577 10824 9608
rect 11149 9605 11161 9608
rect 11195 9636 11207 9639
rect 11195 9608 11652 9636
rect 11195 9605 11207 9608
rect 11149 9599 11207 9605
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 11057 9571 11115 9577
rect 11057 9537 11069 9571
rect 11103 9568 11115 9571
rect 11238 9568 11244 9580
rect 11103 9540 11244 9568
rect 11103 9537 11115 9540
rect 11057 9531 11115 9537
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11624 9577 11652 9608
rect 12268 9577 12296 9646
rect 11609 9571 11667 9577
rect 11609 9537 11621 9571
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 11977 9571 12035 9577
rect 11977 9537 11989 9571
rect 12023 9568 12035 9571
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 12023 9540 12265 9568
rect 12023 9537 12035 9540
rect 11977 9531 12035 9537
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 12434 9534 12440 9586
rect 12492 9574 12498 9586
rect 12492 9568 12572 9574
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12492 9540 12725 9568
rect 12492 9534 12498 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12437 9531 12495 9534
rect 12713 9531 12771 9537
rect 8711 9472 9536 9500
rect 9769 9503 9827 9509
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 9232 9444 9260 9472
rect 9769 9469 9781 9503
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 11701 9503 11759 9509
rect 11701 9469 11713 9503
rect 11747 9500 11759 9503
rect 12066 9500 12072 9512
rect 11747 9472 12072 9500
rect 11747 9469 11759 9472
rect 11701 9463 11759 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 5399 9404 6776 9432
rect 5399 9401 5411 9404
rect 5353 9395 5411 9401
rect 8754 9392 8760 9444
rect 8812 9392 8818 9444
rect 9214 9392 9220 9444
rect 9272 9392 9278 9444
rect 9953 9435 10011 9441
rect 9953 9401 9965 9435
rect 9999 9432 10011 9435
rect 10318 9432 10324 9444
rect 9999 9404 10324 9432
rect 9999 9401 10011 9404
rect 9953 9395 10011 9401
rect 10318 9392 10324 9404
rect 10376 9392 10382 9444
rect 11793 9435 11851 9441
rect 11793 9401 11805 9435
rect 11839 9432 11851 9435
rect 12158 9432 12164 9444
rect 11839 9404 12164 9432
rect 11839 9401 11851 9404
rect 11793 9395 11851 9401
rect 12158 9392 12164 9404
rect 12216 9392 12222 9444
rect 12268 9432 12296 9531
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 12618 9500 12624 9512
rect 12575 9472 12624 9500
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12802 9432 12808 9444
rect 12268 9404 12808 9432
rect 12802 9392 12808 9404
rect 12860 9392 12866 9444
rect 3050 9364 3056 9376
rect 2792 9336 3056 9364
rect 2685 9327 2743 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3326 9324 3332 9376
rect 3384 9364 3390 9376
rect 3789 9367 3847 9373
rect 3789 9364 3801 9367
rect 3384 9336 3801 9364
rect 3384 9324 3390 9336
rect 3789 9333 3801 9336
rect 3835 9333 3847 9367
rect 3789 9327 3847 9333
rect 4522 9324 4528 9376
rect 4580 9364 4586 9376
rect 4706 9364 4712 9376
rect 4580 9336 4712 9364
rect 4580 9324 4586 9336
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 6270 9324 6276 9376
rect 6328 9364 6334 9376
rect 7009 9367 7067 9373
rect 7009 9364 7021 9367
rect 6328 9336 7021 9364
rect 6328 9324 6334 9336
rect 7009 9333 7021 9336
rect 7055 9333 7067 9367
rect 7009 9327 7067 9333
rect 8386 9324 8392 9376
rect 8444 9324 8450 9376
rect 8849 9367 8907 9373
rect 8849 9333 8861 9367
rect 8895 9364 8907 9367
rect 9766 9364 9772 9376
rect 8895 9336 9772 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10962 9324 10968 9376
rect 11020 9364 11026 9376
rect 11885 9367 11943 9373
rect 11885 9364 11897 9367
rect 11020 9336 11897 9364
rect 11020 9324 11026 9336
rect 11885 9333 11897 9336
rect 11931 9333 11943 9367
rect 11885 9327 11943 9333
rect 12621 9367 12679 9373
rect 12621 9333 12633 9367
rect 12667 9364 12679 9367
rect 12710 9364 12716 9376
rect 12667 9336 12716 9364
rect 12667 9333 12679 9336
rect 12621 9327 12679 9333
rect 12710 9324 12716 9336
rect 12768 9324 12774 9376
rect 1104 9274 13340 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 13340 9274
rect 1104 9200 13340 9222
rect 3329 9163 3387 9169
rect 3329 9129 3341 9163
rect 3375 9129 3387 9163
rect 3329 9123 3387 9129
rect 2958 9092 2964 9104
rect 2792 9064 2964 9092
rect 2498 8984 2504 9036
rect 2556 9024 2562 9036
rect 2792 9033 2820 9064
rect 2958 9052 2964 9064
rect 3016 9092 3022 9104
rect 3344 9092 3372 9123
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6822 9160 6828 9172
rect 6144 9132 6828 9160
rect 6144 9120 6150 9132
rect 6822 9120 6828 9132
rect 6880 9120 6886 9172
rect 9398 9120 9404 9172
rect 9456 9120 9462 9172
rect 10962 9120 10968 9172
rect 11020 9160 11026 9172
rect 11333 9163 11391 9169
rect 11333 9160 11345 9163
rect 11020 9132 11345 9160
rect 11020 9120 11026 9132
rect 11333 9129 11345 9132
rect 11379 9129 11391 9163
rect 11333 9123 11391 9129
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 12618 9160 12624 9172
rect 12575 9132 12624 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 12618 9120 12624 9132
rect 12676 9120 12682 9172
rect 12802 9120 12808 9172
rect 12860 9120 12866 9172
rect 3016 9064 3372 9092
rect 6365 9095 6423 9101
rect 3016 9052 3022 9064
rect 6365 9061 6377 9095
rect 6411 9092 6423 9095
rect 7190 9092 7196 9104
rect 6411 9064 7196 9092
rect 6411 9061 6423 9064
rect 6365 9055 6423 9061
rect 7190 9052 7196 9064
rect 7248 9052 7254 9104
rect 2777 9027 2835 9033
rect 2556 8996 2728 9024
rect 2556 8984 2562 8996
rect 2590 8916 2596 8968
rect 2648 8916 2654 8968
rect 2700 8965 2728 8996
rect 2777 8993 2789 9027
rect 2823 8993 2835 9027
rect 2777 8987 2835 8993
rect 2866 8984 2872 9036
rect 2924 8984 2930 9036
rect 8386 9024 8392 9036
rect 6564 8996 8392 9024
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 2961 8959 3019 8965
rect 2961 8925 2973 8959
rect 3007 8956 3019 8959
rect 3602 8956 3608 8968
rect 3007 8928 3608 8956
rect 3007 8925 3019 8928
rect 2961 8919 3019 8925
rect 2608 8888 2636 8916
rect 3528 8897 3556 8928
rect 3602 8916 3608 8928
rect 3660 8956 3666 8968
rect 4614 8956 4620 8968
rect 3660 8928 4620 8956
rect 3660 8916 3666 8928
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4706 8916 4712 8968
rect 4764 8956 4770 8968
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4764 8928 4813 8956
rect 4764 8916 4770 8928
rect 4801 8925 4813 8928
rect 4847 8956 4859 8959
rect 5442 8956 5448 8968
rect 4847 8928 5448 8956
rect 4847 8925 4859 8928
rect 4801 8919 4859 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6270 8916 6276 8968
rect 6328 8916 6334 8968
rect 6564 8965 6592 8996
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 6638 8916 6644 8968
rect 6696 8916 6702 8968
rect 9214 8916 9220 8968
rect 9272 8916 9278 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9858 8956 9864 8968
rect 9447 8928 9864 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9858 8916 9864 8928
rect 9916 8916 9922 8968
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8956 11299 8959
rect 11974 8956 11980 8968
rect 11287 8928 11980 8956
rect 11287 8925 11299 8928
rect 11241 8919 11299 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 12986 8916 12992 8968
rect 13044 8916 13050 8968
rect 3297 8891 3355 8897
rect 3297 8888 3309 8891
rect 2608 8860 3309 8888
rect 3297 8857 3309 8860
rect 3343 8857 3355 8891
rect 3297 8851 3355 8857
rect 3513 8891 3571 8897
rect 3513 8857 3525 8891
rect 3559 8857 3571 8891
rect 3513 8851 3571 8857
rect 4985 8891 5043 8897
rect 4985 8857 4997 8891
rect 5031 8888 5043 8891
rect 5258 8888 5264 8900
rect 5031 8860 5264 8888
rect 5031 8857 5043 8860
rect 4985 8851 5043 8857
rect 5258 8848 5264 8860
rect 5316 8848 5322 8900
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 2280 8792 2513 8820
rect 2280 8780 2286 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 2590 8780 2596 8832
rect 2648 8820 2654 8832
rect 3145 8823 3203 8829
rect 3145 8820 3157 8823
rect 2648 8792 3157 8820
rect 2648 8780 2654 8792
rect 3145 8789 3157 8792
rect 3191 8789 3203 8823
rect 3145 8783 3203 8789
rect 4617 8823 4675 8829
rect 4617 8789 4629 8823
rect 4663 8820 4675 8823
rect 4706 8820 4712 8832
rect 4663 8792 4712 8820
rect 4663 8789 4675 8792
rect 4617 8783 4675 8789
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 6730 8780 6736 8832
rect 6788 8820 6794 8832
rect 6825 8823 6883 8829
rect 6825 8820 6837 8823
rect 6788 8792 6837 8820
rect 6788 8780 6794 8792
rect 6825 8789 6837 8792
rect 6871 8789 6883 8823
rect 6825 8783 6883 8789
rect 1104 8730 13340 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 13340 8730
rect 1104 8656 13340 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2372 8588 3556 8616
rect 2372 8576 2378 8588
rect 2133 8551 2191 8557
rect 2133 8517 2145 8551
rect 2179 8548 2191 8551
rect 2406 8548 2412 8560
rect 2179 8520 2412 8548
rect 2179 8517 2191 8520
rect 2133 8511 2191 8517
rect 2406 8508 2412 8520
rect 2464 8508 2470 8560
rect 2866 8508 2872 8560
rect 2924 8508 2930 8560
rect 3528 8548 3556 8588
rect 3602 8576 3608 8628
rect 3660 8576 3666 8628
rect 4246 8576 4252 8628
rect 4304 8616 4310 8628
rect 4982 8616 4988 8628
rect 4304 8588 4988 8616
rect 4304 8576 4310 8588
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 4264 8548 4292 8576
rect 5905 8551 5963 8557
rect 5905 8548 5917 8551
rect 3528 8520 4292 8548
rect 5474 8520 5917 8548
rect 5905 8517 5917 8520
rect 5951 8517 5963 8551
rect 6546 8548 6552 8560
rect 5905 8511 5963 8517
rect 6012 8520 6552 8548
rect 5534 8440 5540 8492
rect 5592 8480 5598 8492
rect 6012 8489 6040 8520
rect 6546 8508 6552 8520
rect 6604 8548 6610 8560
rect 12345 8551 12403 8557
rect 12345 8548 12357 8551
rect 6604 8520 12357 8548
rect 6604 8508 6610 8520
rect 12345 8517 12357 8520
rect 12391 8548 12403 8551
rect 12391 8520 12756 8548
rect 12391 8517 12403 8520
rect 12345 8511 12403 8517
rect 12728 8492 12756 8520
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5592 8452 6009 8480
rect 5592 8440 5598 8452
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 10318 8440 10324 8492
rect 10376 8480 10382 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 10376 8452 10701 8480
rect 10376 8440 10382 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 12618 8440 12624 8492
rect 12676 8440 12682 8492
rect 12710 8440 12716 8492
rect 12768 8440 12774 8492
rect 1854 8372 1860 8424
rect 1912 8372 1918 8424
rect 3970 8372 3976 8424
rect 4028 8372 4034 8424
rect 4249 8415 4307 8421
rect 4249 8381 4261 8415
rect 4295 8412 4307 8415
rect 4614 8412 4620 8424
rect 4295 8384 4620 8412
rect 4295 8381 4307 8384
rect 4249 8375 4307 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5442 8412 5448 8424
rect 4948 8384 5448 8412
rect 4948 8372 4954 8384
rect 5442 8372 5448 8384
rect 5500 8412 5506 8424
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5500 8384 5733 8412
rect 5500 8372 5506 8384
rect 5721 8381 5733 8384
rect 5767 8381 5779 8415
rect 5721 8375 5779 8381
rect 10597 8415 10655 8421
rect 10597 8381 10609 8415
rect 10643 8412 10655 8415
rect 10962 8412 10968 8424
rect 10643 8384 10968 8412
rect 10643 8381 10655 8384
rect 10597 8375 10655 8381
rect 10962 8372 10968 8384
rect 11020 8372 11026 8424
rect 11054 8372 11060 8424
rect 11112 8412 11118 8424
rect 11149 8415 11207 8421
rect 11149 8412 11161 8415
rect 11112 8384 11161 8412
rect 11112 8372 11118 8384
rect 11149 8381 11161 8384
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 12802 8304 12808 8356
rect 12860 8304 12866 8356
rect 3142 8236 3148 8288
rect 3200 8276 3206 8288
rect 5534 8276 5540 8288
rect 3200 8248 5540 8276
rect 3200 8236 3206 8248
rect 5534 8236 5540 8248
rect 5592 8236 5598 8288
rect 1104 8186 13340 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 13340 8186
rect 1104 8112 13340 8134
rect 2222 8032 2228 8084
rect 2280 8032 2286 8084
rect 2406 8032 2412 8084
rect 2464 8032 2470 8084
rect 2866 8032 2872 8084
rect 2924 8072 2930 8084
rect 2961 8075 3019 8081
rect 2961 8072 2973 8075
rect 2924 8044 2973 8072
rect 2924 8032 2930 8044
rect 2961 8041 2973 8044
rect 3007 8041 3019 8075
rect 2961 8035 3019 8041
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5350 8072 5356 8084
rect 5040 8044 5356 8072
rect 5040 8032 5046 8044
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 7377 8075 7435 8081
rect 7377 8072 7389 8075
rect 6052 8044 7389 8072
rect 6052 8032 6058 8044
rect 7377 8041 7389 8044
rect 7423 8072 7435 8075
rect 7742 8072 7748 8084
rect 7423 8044 7748 8072
rect 7423 8041 7435 8044
rect 7377 8035 7435 8041
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 8021 8075 8079 8081
rect 8021 8041 8033 8075
rect 8067 8072 8079 8075
rect 8665 8075 8723 8081
rect 8665 8072 8677 8075
rect 8067 8044 8677 8072
rect 8067 8041 8079 8044
rect 8021 8035 8079 8041
rect 8665 8041 8677 8044
rect 8711 8041 8723 8075
rect 8665 8035 8723 8041
rect 10410 8032 10416 8084
rect 10468 8072 10474 8084
rect 10505 8075 10563 8081
rect 10505 8072 10517 8075
rect 10468 8044 10517 8072
rect 10468 8032 10474 8044
rect 10505 8041 10517 8044
rect 10551 8041 10563 8075
rect 10505 8035 10563 8041
rect 12066 8032 12072 8084
rect 12124 8072 12130 8084
rect 12529 8075 12587 8081
rect 12529 8072 12541 8075
rect 12124 8044 12541 8072
rect 12124 8032 12130 8044
rect 12529 8041 12541 8044
rect 12575 8041 12587 8075
rect 12529 8035 12587 8041
rect 1854 7964 1860 8016
rect 1912 8004 1918 8016
rect 2774 8004 2780 8016
rect 1912 7976 2780 8004
rect 1912 7964 1918 7976
rect 2774 7964 2780 7976
rect 2832 8004 2838 8016
rect 2832 7976 3556 8004
rect 2832 7964 2838 7976
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 1857 7871 1915 7877
rect 1857 7868 1869 7871
rect 1636 7840 1869 7868
rect 1636 7828 1642 7840
rect 1857 7837 1869 7840
rect 1903 7868 1915 7871
rect 2590 7868 2596 7880
rect 1903 7840 2596 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 2590 7828 2596 7840
rect 2648 7828 2654 7880
rect 2869 7871 2927 7877
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3142 7868 3148 7880
rect 2915 7840 3148 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3528 7877 3556 7976
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 4249 8007 4307 8013
rect 4249 8004 4261 8007
rect 4028 7976 4261 8004
rect 4028 7964 4034 7976
rect 4249 7973 4261 7976
rect 4295 7973 4307 8007
rect 4249 7967 4307 7973
rect 7653 8007 7711 8013
rect 7653 7973 7665 8007
rect 7699 8004 7711 8007
rect 8941 8007 8999 8013
rect 8941 8004 8953 8007
rect 7699 7976 8953 8004
rect 7699 7973 7711 7976
rect 7653 7967 7711 7973
rect 8941 7973 8953 7976
rect 8987 7973 8999 8007
rect 8941 7967 8999 7973
rect 3513 7871 3571 7877
rect 3513 7837 3525 7871
rect 3559 7868 3571 7871
rect 3988 7868 4016 7964
rect 4264 7936 4292 7967
rect 5629 7939 5687 7945
rect 5629 7936 5641 7939
rect 4264 7908 5641 7936
rect 5629 7905 5641 7908
rect 5675 7905 5687 7939
rect 5629 7899 5687 7905
rect 6270 7896 6276 7948
rect 6328 7936 6334 7948
rect 7668 7936 7696 7967
rect 9398 7936 9404 7948
rect 6328 7908 7696 7936
rect 8496 7908 9404 7936
rect 6328 7896 6334 7908
rect 8496 7880 8524 7908
rect 9398 7896 9404 7908
rect 9456 7936 9462 7948
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 9456 7908 9505 7936
rect 9456 7896 9462 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 11054 7896 11060 7948
rect 11112 7896 11118 7948
rect 3559 7840 4016 7868
rect 3559 7837 3571 7840
rect 3513 7831 3571 7837
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 8938 7828 8944 7880
rect 8996 7868 9002 7880
rect 10781 7871 10839 7877
rect 10781 7868 10793 7871
rect 8996 7840 10793 7868
rect 8996 7828 9002 7840
rect 10781 7837 10793 7840
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 12710 7828 12716 7880
rect 12768 7828 12774 7880
rect 4246 7760 4252 7812
rect 4304 7800 4310 7812
rect 4706 7800 4712 7812
rect 4304 7772 4712 7800
rect 4304 7760 4310 7772
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 5537 7803 5595 7809
rect 5537 7769 5549 7803
rect 5583 7769 5595 7803
rect 5537 7763 5595 7769
rect 2225 7735 2283 7741
rect 2225 7701 2237 7735
rect 2271 7732 2283 7735
rect 2682 7732 2688 7744
rect 2271 7704 2688 7732
rect 2271 7701 2283 7704
rect 2225 7695 2283 7701
rect 2682 7692 2688 7704
rect 2740 7692 2746 7744
rect 4430 7692 4436 7744
rect 4488 7732 4494 7744
rect 4890 7732 4896 7744
rect 4488 7704 4896 7732
rect 4488 7692 4494 7704
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5552 7732 5580 7763
rect 5902 7760 5908 7812
rect 5960 7760 5966 7812
rect 6638 7760 6644 7812
rect 6696 7760 6702 7812
rect 8294 7760 8300 7812
rect 8352 7760 8358 7812
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8628 7772 9321 7800
rect 8628 7760 8634 7772
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 10321 7803 10379 7809
rect 10321 7769 10333 7803
rect 10367 7800 10379 7803
rect 11054 7800 11060 7812
rect 10367 7772 11060 7800
rect 10367 7769 10379 7772
rect 10321 7763 10379 7769
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 12805 7803 12863 7809
rect 12805 7800 12817 7803
rect 12282 7772 12817 7800
rect 12805 7769 12817 7772
rect 12851 7769 12863 7803
rect 12805 7763 12863 7769
rect 7282 7732 7288 7744
rect 5552 7704 7288 7732
rect 7282 7692 7288 7704
rect 7340 7692 7346 7744
rect 8021 7735 8079 7741
rect 8021 7701 8033 7735
rect 8067 7732 8079 7735
rect 8110 7732 8116 7744
rect 8067 7704 8116 7732
rect 8067 7701 8079 7704
rect 8021 7695 8079 7701
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8202 7692 8208 7744
rect 8260 7692 8266 7744
rect 8478 7692 8484 7744
rect 8536 7732 8542 7744
rect 9125 7735 9183 7741
rect 9125 7732 9137 7735
rect 8536 7704 9137 7732
rect 8536 7692 8542 7704
rect 9125 7701 9137 7704
rect 9171 7701 9183 7735
rect 9125 7695 9183 7701
rect 9214 7692 9220 7744
rect 9272 7692 9278 7744
rect 10502 7692 10508 7744
rect 10560 7741 10566 7744
rect 10560 7735 10579 7741
rect 10567 7701 10579 7735
rect 10560 7695 10579 7701
rect 10560 7692 10566 7695
rect 10686 7692 10692 7744
rect 10744 7692 10750 7744
rect 1104 7642 13340 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 13340 7642
rect 1104 7568 13340 7590
rect 4433 7531 4491 7537
rect 4433 7497 4445 7531
rect 4479 7528 4491 7531
rect 4522 7528 4528 7540
rect 4479 7500 4528 7528
rect 4479 7497 4491 7500
rect 4433 7491 4491 7497
rect 4522 7488 4528 7500
rect 4580 7488 4586 7540
rect 4693 7531 4751 7537
rect 4693 7497 4705 7531
rect 4739 7528 4751 7531
rect 4739 7500 5856 7528
rect 4739 7497 4751 7500
rect 4693 7491 4751 7497
rect 5828 7472 5856 7500
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 6733 7531 6791 7537
rect 6733 7528 6745 7531
rect 6696 7500 6745 7528
rect 6696 7488 6702 7500
rect 6733 7497 6745 7500
rect 6779 7497 6791 7531
rect 8938 7528 8944 7540
rect 6733 7491 6791 7497
rect 7668 7500 8944 7528
rect 4249 7463 4307 7469
rect 4249 7429 4261 7463
rect 4295 7429 4307 7463
rect 4249 7423 4307 7429
rect 4893 7463 4951 7469
rect 4893 7429 4905 7463
rect 4939 7460 4951 7463
rect 4939 7432 5764 7460
rect 4939 7429 4951 7432
rect 4893 7423 4951 7429
rect 4264 7392 4292 7423
rect 4982 7392 4988 7404
rect 4264 7364 4988 7392
rect 4982 7352 4988 7364
rect 5040 7352 5046 7404
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 5736 7392 5764 7432
rect 5810 7420 5816 7472
rect 5868 7460 5874 7472
rect 6181 7463 6239 7469
rect 6181 7460 6193 7463
rect 5868 7432 6193 7460
rect 5868 7420 5874 7432
rect 6181 7429 6193 7432
rect 6227 7460 6239 7463
rect 6270 7460 6276 7472
rect 6227 7432 6276 7460
rect 6227 7429 6239 7432
rect 6181 7423 6239 7429
rect 6270 7420 6276 7432
rect 6328 7420 6334 7472
rect 5994 7392 6000 7404
rect 5736 7364 6000 7392
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6604 7364 6653 7392
rect 6604 7352 6610 7364
rect 6641 7361 6653 7364
rect 6687 7392 6699 7395
rect 7558 7392 7564 7404
rect 6687 7364 7564 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 7558 7352 7564 7364
rect 7616 7352 7622 7404
rect 7668 7401 7696 7500
rect 8938 7488 8944 7500
rect 8996 7488 9002 7540
rect 9398 7488 9404 7540
rect 9456 7488 9462 7540
rect 11054 7488 11060 7540
rect 11112 7488 11118 7540
rect 11146 7488 11152 7540
rect 11204 7528 11210 7540
rect 11204 7500 11744 7528
rect 11204 7488 11210 7500
rect 7929 7463 7987 7469
rect 7929 7429 7941 7463
rect 7975 7460 7987 7463
rect 8202 7460 8208 7472
rect 7975 7432 8208 7460
rect 7975 7429 7987 7432
rect 7929 7423 7987 7429
rect 8202 7420 8208 7432
rect 8260 7420 8266 7472
rect 9585 7463 9643 7469
rect 9585 7460 9597 7463
rect 9154 7432 9597 7460
rect 9585 7429 9597 7432
rect 9631 7429 9643 7463
rect 9585 7423 9643 7429
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 11716 7469 11744 7500
rect 11517 7463 11575 7469
rect 11517 7460 11529 7463
rect 10560 7432 11529 7460
rect 10560 7420 10566 7432
rect 11517 7429 11529 7432
rect 11563 7429 11575 7463
rect 11517 7423 11575 7429
rect 11701 7463 11759 7469
rect 11701 7429 11713 7463
rect 11747 7460 11759 7463
rect 11974 7460 11980 7472
rect 11747 7432 11980 7460
rect 11747 7429 11759 7432
rect 11701 7423 11759 7429
rect 11974 7420 11980 7432
rect 12032 7420 12038 7472
rect 7653 7395 7711 7401
rect 7653 7361 7665 7395
rect 7699 7361 7711 7395
rect 7653 7355 7711 7361
rect 9674 7352 9680 7404
rect 9732 7352 9738 7404
rect 11057 7395 11115 7401
rect 11057 7361 11069 7395
rect 11103 7392 11115 7395
rect 11146 7392 11152 7404
rect 11103 7364 11152 7392
rect 11103 7361 11115 7364
rect 11057 7355 11115 7361
rect 11146 7352 11152 7364
rect 11204 7352 11210 7404
rect 11238 7352 11244 7404
rect 11296 7401 11302 7404
rect 11296 7395 11309 7401
rect 11297 7392 11309 7395
rect 11885 7395 11943 7401
rect 11885 7392 11897 7395
rect 11297 7364 11897 7392
rect 11297 7361 11309 7364
rect 11296 7355 11309 7361
rect 11885 7361 11897 7364
rect 11931 7392 11943 7395
rect 12066 7392 12072 7404
rect 11931 7364 12072 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 11296 7352 11302 7355
rect 12066 7352 12072 7364
rect 12124 7352 12130 7404
rect 5350 7284 5356 7336
rect 5408 7324 5414 7336
rect 10318 7324 10324 7336
rect 5408 7296 10324 7324
rect 5408 7284 5414 7296
rect 9048 7268 9076 7296
rect 10318 7284 10324 7296
rect 10376 7284 10382 7336
rect 12526 7284 12532 7336
rect 12584 7284 12590 7336
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 4525 7259 4583 7265
rect 4525 7256 4537 7259
rect 3936 7228 4537 7256
rect 3936 7216 3942 7228
rect 4525 7225 4537 7228
rect 4571 7225 4583 7259
rect 4525 7219 4583 7225
rect 9030 7216 9036 7268
rect 9088 7216 9094 7268
rect 4246 7148 4252 7200
rect 4304 7148 4310 7200
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 4709 7191 4767 7197
rect 4709 7188 4721 7191
rect 4672 7160 4721 7188
rect 4672 7148 4678 7160
rect 4709 7157 4721 7160
rect 4755 7157 4767 7191
rect 4709 7151 4767 7157
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 5813 7191 5871 7197
rect 5813 7188 5825 7191
rect 5408 7160 5825 7188
rect 5408 7148 5414 7160
rect 5813 7157 5825 7160
rect 5859 7157 5871 7191
rect 5813 7151 5871 7157
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12069 7191 12127 7197
rect 12069 7188 12081 7191
rect 12032 7160 12081 7188
rect 12032 7148 12038 7160
rect 12069 7157 12081 7160
rect 12115 7157 12127 7191
rect 12069 7151 12127 7157
rect 1104 7098 13340 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 13340 7098
rect 1104 7024 13340 7046
rect 5350 6944 5356 6996
rect 5408 6944 5414 6996
rect 5537 6987 5595 6993
rect 5537 6953 5549 6987
rect 5583 6984 5595 6987
rect 5902 6984 5908 6996
rect 5583 6956 5908 6984
rect 5583 6953 5595 6956
rect 5537 6947 5595 6953
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7745 6987 7803 6993
rect 7745 6984 7757 6987
rect 7340 6956 7757 6984
rect 7340 6944 7346 6956
rect 7745 6953 7757 6956
rect 7791 6984 7803 6987
rect 8202 6984 8208 6996
rect 7791 6956 8208 6984
rect 7791 6953 7803 6956
rect 7745 6947 7803 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8294 6944 8300 6996
rect 8352 6944 8358 6996
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6984 8539 6987
rect 9214 6984 9220 6996
rect 8527 6956 9220 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 9214 6944 9220 6956
rect 9272 6984 9278 6996
rect 9398 6984 9404 6996
rect 9272 6956 9404 6984
rect 9272 6944 9278 6956
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 10686 6944 10692 6996
rect 10744 6984 10750 6996
rect 11314 6987 11372 6993
rect 11314 6984 11326 6987
rect 10744 6956 11326 6984
rect 10744 6944 10750 6956
rect 11314 6953 11326 6956
rect 11360 6953 11372 6987
rect 11314 6947 11372 6953
rect 12526 6944 12532 6996
rect 12584 6984 12590 6996
rect 12805 6987 12863 6993
rect 12805 6984 12817 6987
rect 12584 6956 12817 6984
rect 12584 6944 12590 6956
rect 12805 6953 12817 6956
rect 12851 6953 12863 6987
rect 12805 6947 12863 6953
rect 4982 6916 4988 6928
rect 4724 6888 4988 6916
rect 2682 6808 2688 6860
rect 2740 6848 2746 6860
rect 4724 6848 4752 6888
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 6089 6919 6147 6925
rect 6089 6885 6101 6919
rect 6135 6885 6147 6919
rect 6089 6879 6147 6885
rect 2740 6820 4752 6848
rect 4801 6851 4859 6857
rect 2740 6808 2746 6820
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 6104 6848 6132 6879
rect 4847 6820 6132 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 8938 6808 8944 6860
rect 8996 6848 9002 6860
rect 11057 6851 11115 6857
rect 11057 6848 11069 6851
rect 8996 6820 11069 6848
rect 8996 6808 9002 6820
rect 11057 6817 11069 6820
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1578 6740 1584 6792
rect 1636 6780 1642 6792
rect 2133 6783 2191 6789
rect 2133 6780 2145 6783
rect 1636 6752 2145 6780
rect 1636 6740 1642 6752
rect 2133 6749 2145 6752
rect 2179 6780 2191 6783
rect 2590 6780 2596 6792
rect 2179 6752 2596 6780
rect 2179 6749 2191 6752
rect 2133 6743 2191 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 3142 6780 3148 6792
rect 2915 6752 3148 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 4706 6740 4712 6792
rect 4764 6740 4770 6792
rect 4985 6783 5043 6789
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5258 6780 5264 6792
rect 5031 6752 5264 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5258 6740 5264 6752
rect 5316 6780 5322 6792
rect 5629 6783 5687 6789
rect 5629 6780 5641 6783
rect 5316 6752 5641 6780
rect 5316 6740 5322 6752
rect 5629 6749 5641 6752
rect 5675 6749 5687 6783
rect 5629 6743 5687 6749
rect 5810 6740 5816 6792
rect 5868 6740 5874 6792
rect 5994 6740 6000 6792
rect 6052 6740 6058 6792
rect 6178 6740 6184 6792
rect 6236 6780 6242 6792
rect 6273 6783 6331 6789
rect 6273 6780 6285 6783
rect 6236 6752 6285 6780
rect 6236 6740 6242 6752
rect 6273 6749 6285 6752
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6454 6740 6460 6792
rect 6512 6740 6518 6792
rect 1486 6672 1492 6724
rect 1544 6712 1550 6724
rect 2317 6715 2375 6721
rect 2317 6712 2329 6715
rect 1544 6684 2329 6712
rect 1544 6672 1550 6684
rect 2317 6681 2329 6684
rect 2363 6681 2375 6715
rect 4798 6712 4804 6724
rect 2317 6675 2375 6681
rect 2424 6684 4804 6712
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2424 6644 2452 6684
rect 4798 6672 4804 6684
rect 4856 6672 4862 6724
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 6196 6712 6224 6740
rect 8478 6721 8484 6724
rect 5776 6684 6224 6712
rect 8465 6715 8484 6721
rect 5776 6672 5782 6684
rect 8465 6681 8477 6715
rect 8465 6675 8484 6681
rect 8478 6672 8484 6675
rect 8536 6672 8542 6724
rect 8570 6672 8576 6724
rect 8628 6712 8634 6724
rect 8665 6715 8723 6721
rect 8665 6712 8677 6715
rect 8628 6684 8677 6712
rect 8628 6672 8634 6684
rect 8665 6681 8677 6684
rect 8711 6681 8723 6715
rect 8665 6675 8723 6681
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 9217 6715 9275 6721
rect 9217 6712 9229 6715
rect 8812 6684 9229 6712
rect 8812 6672 8818 6684
rect 9217 6681 9229 6684
rect 9263 6681 9275 6715
rect 12802 6712 12808 6724
rect 9217 6675 9275 6681
rect 9324 6684 9706 6712
rect 12558 6684 12808 6712
rect 1627 6616 2452 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 2961 6647 3019 6653
rect 2961 6644 2973 6647
rect 2924 6616 2973 6644
rect 2924 6604 2930 6616
rect 2961 6613 2973 6616
rect 3007 6613 3019 6647
rect 2961 6607 3019 6613
rect 4338 6604 4344 6656
rect 4396 6604 4402 6656
rect 4982 6604 4988 6656
rect 5040 6644 5046 6656
rect 5353 6647 5411 6653
rect 5353 6644 5365 6647
rect 5040 6616 5365 6644
rect 5040 6604 5046 6616
rect 5353 6613 5365 6616
rect 5399 6644 5411 6647
rect 7926 6644 7932 6656
rect 5399 6616 7932 6644
rect 5399 6613 5411 6616
rect 5353 6607 5411 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8846 6604 8852 6656
rect 8904 6644 8910 6656
rect 9324 6644 9352 6684
rect 12802 6672 12808 6684
rect 12860 6672 12866 6724
rect 8904 6616 9352 6644
rect 8904 6604 8910 6616
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 9456 6616 10701 6644
rect 9456 6604 9462 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 1104 6554 13340 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 13340 6554
rect 1104 6480 13340 6502
rect 1486 6400 1492 6452
rect 1544 6440 1550 6452
rect 1544 6412 3648 6440
rect 1544 6400 1550 6412
rect 2866 6332 2872 6384
rect 2924 6332 2930 6384
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 1854 6264 1860 6316
rect 1912 6264 1918 6316
rect 2130 6196 2136 6248
rect 2188 6196 2194 6248
rect 3620 6177 3648 6412
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5721 6443 5779 6449
rect 5721 6440 5733 6443
rect 4764 6412 5733 6440
rect 4764 6400 4770 6412
rect 5721 6409 5733 6412
rect 5767 6409 5779 6443
rect 5721 6403 5779 6409
rect 6733 6443 6791 6449
rect 6733 6409 6745 6443
rect 6779 6440 6791 6443
rect 6822 6440 6828 6452
rect 6779 6412 6828 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8754 6440 8760 6452
rect 8343 6412 8760 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8754 6400 8760 6412
rect 8812 6400 8818 6452
rect 8938 6400 8944 6452
rect 8996 6440 9002 6452
rect 9582 6440 9588 6452
rect 8996 6412 9588 6440
rect 8996 6400 9002 6412
rect 9582 6400 9588 6412
rect 9640 6440 9646 6452
rect 9677 6443 9735 6449
rect 9677 6440 9689 6443
rect 9640 6412 9689 6440
rect 9640 6400 9646 6412
rect 9677 6409 9689 6412
rect 9723 6409 9735 6443
rect 9677 6403 9735 6409
rect 10226 6400 10232 6452
rect 10284 6440 10290 6452
rect 10387 6443 10445 6449
rect 10387 6440 10399 6443
rect 10284 6412 10399 6440
rect 10284 6400 10290 6412
rect 10387 6409 10399 6412
rect 10433 6440 10445 6443
rect 10965 6443 11023 6449
rect 10965 6440 10977 6443
rect 10433 6412 10977 6440
rect 10433 6409 10445 6412
rect 10387 6403 10445 6409
rect 10965 6409 10977 6412
rect 11011 6440 11023 6443
rect 11146 6440 11152 6452
rect 11011 6412 11152 6440
rect 11011 6409 11023 6412
rect 10965 6403 11023 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 4798 6332 4804 6384
rect 4856 6372 4862 6384
rect 4856 6344 5580 6372
rect 4856 6332 4862 6344
rect 4338 6264 4344 6316
rect 4396 6304 4402 6316
rect 4614 6304 4620 6316
rect 4396 6276 4620 6304
rect 4396 6264 4402 6276
rect 4614 6264 4620 6276
rect 4672 6304 4678 6316
rect 5552 6313 5580 6344
rect 8110 6332 8116 6384
rect 8168 6332 8174 6384
rect 8202 6332 8208 6384
rect 8260 6372 8266 6384
rect 8389 6375 8447 6381
rect 8389 6372 8401 6375
rect 8260 6344 8401 6372
rect 8260 6332 8266 6344
rect 8389 6341 8401 6344
rect 8435 6341 8447 6375
rect 8389 6335 8447 6341
rect 10597 6375 10655 6381
rect 10597 6341 10609 6375
rect 10643 6372 10655 6375
rect 11238 6372 11244 6384
rect 10643 6344 11244 6372
rect 10643 6341 10655 6344
rect 10597 6335 10655 6341
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 12066 6332 12072 6384
rect 12124 6332 12130 6384
rect 4985 6307 5043 6313
rect 4985 6304 4997 6307
rect 4672 6276 4997 6304
rect 4672 6264 4678 6276
rect 4985 6273 4997 6276
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 5537 6307 5595 6313
rect 5537 6273 5549 6307
rect 5583 6304 5595 6307
rect 5629 6307 5687 6313
rect 5629 6304 5641 6307
rect 5583 6276 5641 6304
rect 5583 6273 5595 6276
rect 5537 6267 5595 6273
rect 5629 6273 5641 6276
rect 5675 6273 5687 6307
rect 5629 6267 5687 6273
rect 5905 6307 5963 6313
rect 5905 6273 5917 6307
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 4801 6239 4859 6245
rect 4801 6205 4813 6239
rect 4847 6205 4859 6239
rect 4801 6199 4859 6205
rect 3605 6171 3663 6177
rect 3605 6137 3617 6171
rect 3651 6168 3663 6171
rect 3970 6168 3976 6180
rect 3651 6140 3976 6168
rect 3651 6137 3663 6140
rect 3605 6131 3663 6137
rect 3970 6128 3976 6140
rect 4028 6168 4034 6180
rect 4816 6168 4844 6199
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 5261 6239 5319 6245
rect 5261 6236 5273 6239
rect 5132 6208 5273 6236
rect 5132 6196 5138 6208
rect 5261 6205 5273 6208
rect 5307 6236 5319 6239
rect 5442 6236 5448 6248
rect 5307 6208 5448 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5920 6168 5948 6267
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6546 6313 6552 6316
rect 6519 6307 6552 6313
rect 6519 6273 6531 6307
rect 6519 6267 6552 6273
rect 6546 6264 6552 6267
rect 6604 6264 6610 6316
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 7745 6307 7803 6313
rect 7745 6273 7757 6307
rect 7791 6304 7803 6307
rect 8294 6304 8300 6316
rect 7791 6276 8300 6304
rect 7791 6273 7803 6276
rect 7745 6267 7803 6273
rect 8294 6264 8300 6276
rect 8352 6264 8358 6316
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9674 6304 9680 6316
rect 8628 6276 9680 6304
rect 8628 6264 8634 6276
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 10870 6264 10876 6316
rect 10928 6264 10934 6316
rect 11057 6307 11115 6313
rect 11057 6273 11069 6307
rect 11103 6304 11115 6307
rect 12526 6304 12532 6316
rect 11103 6276 12532 6304
rect 11103 6273 11115 6276
rect 11057 6267 11115 6273
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 10689 6239 10747 6245
rect 10689 6236 10701 6239
rect 9548 6208 10701 6236
rect 9548 6196 9554 6208
rect 10689 6205 10701 6208
rect 10735 6205 10747 6239
rect 10689 6199 10747 6205
rect 11072 6168 11100 6267
rect 12526 6264 12532 6276
rect 12584 6304 12590 6316
rect 12621 6307 12679 6313
rect 12621 6304 12633 6307
rect 12584 6276 12633 6304
rect 12584 6264 12590 6276
rect 12621 6273 12633 6276
rect 12667 6273 12679 6307
rect 12621 6267 12679 6273
rect 4028 6140 5948 6168
rect 10428 6140 11100 6168
rect 4028 6128 4034 6140
rect 1765 6103 1823 6109
rect 1765 6069 1777 6103
rect 1811 6100 1823 6103
rect 2866 6100 2872 6112
rect 1811 6072 2872 6100
rect 1811 6069 1823 6072
rect 1765 6063 1823 6069
rect 2866 6060 2872 6072
rect 2924 6060 2930 6112
rect 5169 6103 5227 6109
rect 5169 6069 5181 6103
rect 5215 6100 5227 6103
rect 5258 6100 5264 6112
rect 5215 6072 5264 6100
rect 5215 6069 5227 6072
rect 5169 6063 5227 6069
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5350 6060 5356 6112
rect 5408 6060 5414 6112
rect 5445 6103 5503 6109
rect 5445 6069 5457 6103
rect 5491 6100 5503 6103
rect 5718 6100 5724 6112
rect 5491 6072 5724 6100
rect 5491 6069 5503 6072
rect 5445 6063 5503 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5994 6060 6000 6112
rect 6052 6060 6058 6112
rect 6917 6103 6975 6109
rect 6917 6069 6929 6103
rect 6963 6100 6975 6103
rect 7006 6100 7012 6112
rect 6963 6072 7012 6100
rect 6963 6069 6975 6072
rect 6917 6063 6975 6069
rect 7006 6060 7012 6072
rect 7064 6060 7070 6112
rect 8113 6103 8171 6109
rect 8113 6069 8125 6103
rect 8159 6100 8171 6103
rect 8938 6100 8944 6112
rect 8159 6072 8944 6100
rect 8159 6069 8171 6072
rect 8113 6063 8171 6069
rect 8938 6060 8944 6072
rect 8996 6060 9002 6112
rect 10226 6060 10232 6112
rect 10284 6060 10290 6112
rect 10428 6109 10456 6140
rect 10413 6103 10471 6109
rect 10413 6069 10425 6103
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 11698 6100 11704 6112
rect 10928 6072 11704 6100
rect 10928 6060 10934 6072
rect 11698 6060 11704 6072
rect 11756 6060 11762 6112
rect 1104 6010 13340 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 13340 6010
rect 1104 5936 13340 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 2188 5868 2329 5896
rect 2188 5856 2194 5868
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 2317 5859 2375 5865
rect 2498 5856 2504 5908
rect 2556 5856 2562 5908
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 6454 5896 6460 5908
rect 5092 5868 6460 5896
rect 2866 5788 2872 5840
rect 2924 5788 2930 5840
rect 4798 5788 4804 5840
rect 4856 5828 4862 5840
rect 4893 5831 4951 5837
rect 4893 5828 4905 5831
rect 4856 5800 4905 5828
rect 4856 5788 4862 5800
rect 4893 5797 4905 5800
rect 4939 5797 4951 5831
rect 4893 5791 4951 5797
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5692 2191 5695
rect 2774 5692 2780 5704
rect 2179 5664 2780 5692
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2774 5652 2780 5664
rect 2832 5652 2838 5704
rect 2884 5692 2912 5788
rect 2961 5695 3019 5701
rect 2961 5692 2973 5695
rect 2884 5664 2973 5692
rect 2961 5661 2973 5664
rect 3007 5661 3019 5695
rect 2961 5655 3019 5661
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5692 3203 5695
rect 3191 5664 4200 5692
rect 3191 5661 3203 5664
rect 3145 5655 3203 5661
rect 4172 5636 4200 5664
rect 4706 5652 4712 5704
rect 4764 5652 4770 5704
rect 5092 5701 5120 5868
rect 6454 5856 6460 5868
rect 6512 5856 6518 5908
rect 6546 5856 6552 5908
rect 6604 5856 6610 5908
rect 7190 5856 7196 5908
rect 7248 5896 7254 5908
rect 7285 5899 7343 5905
rect 7285 5896 7297 5899
rect 7248 5868 7297 5896
rect 7248 5856 7254 5868
rect 7285 5865 7297 5868
rect 7331 5865 7343 5899
rect 7285 5859 7343 5865
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5896 8723 5899
rect 8846 5896 8852 5908
rect 8711 5868 8852 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 8846 5856 8852 5868
rect 8904 5856 8910 5908
rect 8938 5856 8944 5908
rect 8996 5856 9002 5908
rect 9950 5856 9956 5908
rect 10008 5856 10014 5908
rect 10413 5899 10471 5905
rect 10413 5865 10425 5899
rect 10459 5896 10471 5899
rect 11514 5896 11520 5908
rect 10459 5868 11520 5896
rect 10459 5865 10471 5868
rect 10413 5859 10471 5865
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 12621 5899 12679 5905
rect 12621 5896 12633 5899
rect 11756 5868 12633 5896
rect 11756 5856 11762 5868
rect 12621 5865 12633 5868
rect 12667 5865 12679 5899
rect 12621 5859 12679 5865
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 5224 5800 5396 5828
rect 5224 5788 5230 5800
rect 4985 5695 5043 5701
rect 4985 5694 4997 5695
rect 4816 5666 4997 5694
rect 1765 5627 1823 5633
rect 1765 5593 1777 5627
rect 1811 5624 1823 5627
rect 2501 5627 2559 5633
rect 2501 5624 2513 5627
rect 1811 5596 2513 5624
rect 1811 5593 1823 5596
rect 1765 5587 1823 5593
rect 2501 5593 2513 5596
rect 2547 5624 2559 5627
rect 2682 5624 2688 5636
rect 2547 5596 2688 5624
rect 2547 5593 2559 5596
rect 2501 5587 2559 5593
rect 2682 5584 2688 5596
rect 2740 5584 2746 5636
rect 3941 5627 3999 5633
rect 3941 5624 3953 5627
rect 3252 5596 3953 5624
rect 2590 5516 2596 5568
rect 2648 5556 2654 5568
rect 3252 5556 3280 5596
rect 3941 5593 3953 5596
rect 3987 5593 3999 5627
rect 3941 5587 3999 5593
rect 4154 5584 4160 5636
rect 4212 5584 4218 5636
rect 4816 5624 4844 5666
rect 4985 5661 4997 5666
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5166 5652 5172 5704
rect 5224 5692 5230 5704
rect 5368 5701 5396 5800
rect 5442 5788 5448 5840
rect 5500 5828 5506 5840
rect 6086 5828 6092 5840
rect 5500 5800 6092 5828
rect 5500 5788 5506 5800
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 7006 5828 7012 5840
rect 6196 5800 7012 5828
rect 6196 5769 6224 5800
rect 7006 5788 7012 5800
rect 7064 5788 7070 5840
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 9306 5828 9312 5840
rect 8536 5800 9312 5828
rect 8536 5788 8542 5800
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 9582 5788 9588 5840
rect 9640 5788 9646 5840
rect 10226 5788 10232 5840
rect 10284 5828 10290 5840
rect 10781 5831 10839 5837
rect 10781 5828 10793 5831
rect 10284 5800 10793 5828
rect 10284 5788 10290 5800
rect 10781 5797 10793 5800
rect 10827 5828 10839 5831
rect 10827 5800 11008 5828
rect 10827 5797 10839 5800
rect 10781 5791 10839 5797
rect 6181 5763 6239 5769
rect 6181 5760 6193 5763
rect 5736 5732 6193 5760
rect 5353 5695 5411 5701
rect 5224 5664 5269 5692
rect 5224 5652 5230 5664
rect 5353 5661 5365 5695
rect 5399 5661 5411 5695
rect 5353 5655 5411 5661
rect 5581 5695 5639 5701
rect 5581 5661 5593 5695
rect 5627 5686 5639 5695
rect 5736 5686 5764 5732
rect 6181 5729 6193 5732
rect 6227 5729 6239 5763
rect 6181 5723 6239 5729
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6917 5763 6975 5769
rect 6917 5760 6929 5763
rect 6512 5732 6929 5760
rect 6512 5720 6518 5732
rect 6917 5729 6929 5732
rect 6963 5729 6975 5763
rect 9600 5760 9628 5788
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 6917 5723 6975 5729
rect 8404 5732 9444 5760
rect 9600 5732 10885 5760
rect 8404 5704 8432 5732
rect 5627 5661 5764 5686
rect 5581 5658 5764 5661
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5661 5871 5695
rect 5581 5655 5639 5658
rect 5813 5655 5871 5661
rect 5184 5624 5212 5652
rect 4816 5596 5212 5624
rect 5445 5627 5503 5633
rect 5445 5593 5457 5627
rect 5491 5624 5503 5627
rect 5828 5624 5856 5655
rect 5994 5652 6000 5704
rect 6052 5652 6058 5704
rect 6086 5652 6092 5704
rect 6144 5652 6150 5704
rect 6365 5695 6423 5701
rect 6365 5661 6377 5695
rect 6411 5692 6423 5695
rect 6546 5692 6552 5704
rect 6411 5664 6552 5692
rect 6411 5661 6423 5664
rect 6365 5655 6423 5661
rect 6546 5652 6552 5664
rect 6604 5652 6610 5704
rect 6638 5652 6644 5704
rect 6696 5652 6702 5704
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7190 5692 7196 5704
rect 7147 5664 7196 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 6656 5624 6684 5652
rect 5491 5596 5672 5624
rect 5828 5596 6684 5624
rect 5491 5593 5503 5596
rect 5445 5587 5503 5593
rect 5644 5568 5672 5596
rect 2648 5528 3280 5556
rect 2648 5516 2654 5528
rect 3326 5516 3332 5568
rect 3384 5516 3390 5568
rect 3694 5516 3700 5568
rect 3752 5556 3758 5568
rect 3789 5559 3847 5565
rect 3789 5556 3801 5559
rect 3752 5528 3801 5556
rect 3752 5516 3758 5528
rect 3789 5525 3801 5528
rect 3835 5525 3847 5559
rect 3789 5519 3847 5525
rect 4338 5516 4344 5568
rect 4396 5556 4402 5568
rect 4525 5559 4583 5565
rect 4525 5556 4537 5559
rect 4396 5528 4537 5556
rect 4396 5516 4402 5528
rect 4525 5525 4537 5528
rect 4571 5556 4583 5559
rect 4798 5556 4804 5568
rect 4571 5528 4804 5556
rect 4571 5525 4583 5528
rect 4525 5519 4583 5525
rect 4798 5516 4804 5528
rect 4856 5556 4862 5568
rect 5534 5556 5540 5568
rect 4856 5528 5540 5556
rect 4856 5516 4862 5528
rect 5534 5516 5540 5528
rect 5592 5516 5598 5568
rect 5626 5516 5632 5568
rect 5684 5516 5690 5568
rect 5721 5559 5779 5565
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 6362 5556 6368 5568
rect 5767 5528 6368 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 6362 5516 6368 5528
rect 6420 5556 6426 5568
rect 6840 5556 6868 5655
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5692 8355 5695
rect 8386 5692 8392 5704
rect 8343 5664 8392 5692
rect 8343 5661 8355 5664
rect 8297 5655 8355 5661
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8478 5652 8484 5704
rect 8536 5652 8542 5704
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 9125 5695 9183 5701
rect 9125 5661 9137 5695
rect 9171 5692 9183 5695
rect 9214 5692 9220 5704
rect 9171 5664 9220 5692
rect 9171 5661 9183 5664
rect 9125 5655 9183 5661
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 9416 5701 9444 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 10980 5760 11008 5800
rect 11238 5760 11244 5772
rect 10980 5732 11244 5760
rect 10873 5723 10931 5729
rect 11238 5720 11244 5732
rect 11296 5720 11302 5772
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5692 9459 5695
rect 9490 5692 9496 5704
rect 9447 5664 9496 5692
rect 9447 5661 9459 5664
rect 9401 5655 9459 5661
rect 9490 5652 9496 5664
rect 9548 5692 9554 5704
rect 9585 5695 9643 5701
rect 9585 5692 9597 5695
rect 9548 5664 9597 5692
rect 9548 5652 9554 5664
rect 9585 5661 9597 5664
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 8110 5584 8116 5636
rect 8168 5624 8174 5636
rect 8662 5624 8668 5636
rect 8168 5596 8668 5624
rect 8168 5584 8174 5596
rect 8662 5584 8668 5596
rect 8720 5624 8726 5636
rect 9953 5627 10011 5633
rect 9953 5624 9965 5627
rect 8720 5596 9965 5624
rect 8720 5584 8726 5596
rect 9416 5568 9444 5596
rect 9953 5593 9965 5596
rect 9999 5624 10011 5627
rect 10042 5624 10048 5636
rect 9999 5596 10048 5624
rect 9999 5593 10011 5596
rect 9953 5587 10011 5593
rect 10042 5584 10048 5596
rect 10100 5584 10106 5636
rect 10778 5624 10784 5636
rect 10152 5596 10784 5624
rect 6420 5528 6868 5556
rect 6420 5516 6426 5528
rect 8478 5516 8484 5568
rect 8536 5516 8542 5568
rect 9306 5516 9312 5568
rect 9364 5516 9370 5568
rect 9398 5516 9404 5568
rect 9456 5516 9462 5568
rect 10152 5565 10180 5596
rect 10778 5584 10784 5596
rect 10836 5584 10842 5636
rect 11054 5584 11060 5636
rect 11112 5624 11118 5636
rect 11149 5627 11207 5633
rect 11149 5624 11161 5627
rect 11112 5596 11161 5624
rect 11112 5584 11118 5596
rect 11149 5593 11161 5596
rect 11195 5593 11207 5627
rect 12802 5624 12808 5636
rect 12374 5596 12808 5624
rect 11149 5587 11207 5593
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 10137 5559 10195 5565
rect 10137 5525 10149 5559
rect 10183 5525 10195 5559
rect 10137 5519 10195 5525
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 10410 5516 10416 5568
rect 10468 5516 10474 5568
rect 1104 5466 13340 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 13340 5466
rect 1104 5392 13340 5414
rect 4614 5352 4620 5364
rect 4080 5324 4620 5352
rect 3786 5284 3792 5296
rect 3358 5256 3792 5284
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 4080 5284 4108 5324
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 4706 5312 4712 5364
rect 4764 5352 4770 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 4764 5324 4813 5352
rect 4764 5312 4770 5324
rect 4801 5321 4813 5324
rect 4847 5321 4859 5355
rect 4801 5315 4859 5321
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 5350 5352 5356 5364
rect 4948 5324 5356 5352
rect 4948 5312 4954 5324
rect 5350 5312 5356 5324
rect 5408 5352 5414 5364
rect 5971 5355 6029 5361
rect 5971 5352 5983 5355
rect 5408 5324 5983 5352
rect 5408 5312 5414 5324
rect 5971 5321 5983 5324
rect 6017 5321 6029 5355
rect 5971 5315 6029 5321
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 7190 5352 7196 5364
rect 6604 5324 7196 5352
rect 6604 5312 6610 5324
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 11514 5312 11520 5364
rect 11572 5312 11578 5364
rect 12802 5312 12808 5364
rect 12860 5312 12866 5364
rect 3988 5256 4108 5284
rect 4249 5287 4307 5293
rect 1854 5176 1860 5228
rect 1912 5176 1918 5228
rect 3988 5225 4016 5256
rect 4249 5253 4261 5287
rect 4295 5284 4307 5287
rect 4985 5287 5043 5293
rect 4985 5284 4997 5287
rect 4295 5256 4997 5284
rect 4295 5253 4307 5256
rect 4249 5247 4307 5253
rect 4985 5253 4997 5256
rect 5031 5284 5043 5287
rect 5031 5256 5442 5284
rect 5031 5253 5043 5256
rect 4985 5247 5043 5253
rect 5414 5238 5442 5256
rect 5626 5244 5632 5296
rect 5684 5284 5690 5296
rect 6181 5287 6239 5293
rect 6181 5284 6193 5287
rect 5684 5256 6193 5284
rect 5684 5244 5690 5256
rect 6181 5253 6193 5256
rect 6227 5253 6239 5287
rect 6181 5247 6239 5253
rect 8662 5244 8668 5296
rect 8720 5244 8726 5296
rect 8881 5287 8939 5293
rect 8881 5253 8893 5287
rect 8927 5284 8939 5287
rect 9125 5287 9183 5293
rect 9125 5284 9137 5287
rect 8927 5256 9137 5284
rect 8927 5253 8939 5256
rect 8881 5247 8939 5253
rect 9125 5253 9137 5256
rect 9171 5253 9183 5287
rect 9125 5247 9183 5253
rect 9490 5244 9496 5296
rect 9548 5244 9554 5296
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 11885 5287 11943 5293
rect 11885 5284 11897 5287
rect 11388 5256 11897 5284
rect 11388 5244 11394 5256
rect 11885 5253 11897 5256
rect 11931 5253 11943 5287
rect 11885 5247 11943 5253
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 3881 5219 3939 5225
rect 3881 5185 3893 5219
rect 3927 5216 3939 5219
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3927 5188 3985 5216
rect 3927 5185 3939 5188
rect 3881 5179 3939 5185
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 2130 5108 2136 5160
rect 2188 5108 2194 5160
rect 3712 5148 3740 5179
rect 4062 5176 4068 5228
rect 4120 5176 4126 5228
rect 4338 5176 4344 5228
rect 4396 5176 4402 5228
rect 5414 5216 5534 5238
rect 5414 5210 5856 5216
rect 5506 5188 5856 5210
rect 4080 5148 4108 5176
rect 5353 5151 5411 5157
rect 5353 5148 5365 5151
rect 3712 5120 4108 5148
rect 4632 5120 5365 5148
rect 3881 5083 3939 5089
rect 3881 5049 3893 5083
rect 3927 5080 3939 5083
rect 4632 5080 4660 5120
rect 5353 5117 5365 5120
rect 5399 5117 5411 5151
rect 5353 5111 5411 5117
rect 3927 5052 4660 5080
rect 3927 5049 3939 5052
rect 3881 5043 3939 5049
rect 5258 5040 5264 5092
rect 5316 5040 5322 5092
rect 5828 5089 5856 5188
rect 9306 5176 9312 5228
rect 9364 5176 9370 5228
rect 9582 5176 9588 5228
rect 9640 5176 9646 5228
rect 10962 5176 10968 5228
rect 11020 5176 11026 5228
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 9861 5151 9919 5157
rect 9861 5117 9873 5151
rect 9907 5148 9919 5151
rect 10226 5148 10232 5160
rect 9907 5120 10232 5148
rect 9907 5117 9919 5120
rect 9861 5111 9919 5117
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 11146 5108 11152 5160
rect 11204 5148 11210 5160
rect 11333 5151 11391 5157
rect 11333 5148 11345 5151
rect 11204 5120 11345 5148
rect 11204 5108 11210 5120
rect 11333 5117 11345 5120
rect 11379 5148 11391 5151
rect 11716 5148 11744 5179
rect 11974 5176 11980 5228
rect 12032 5176 12038 5228
rect 12253 5219 12311 5225
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12618 5216 12624 5228
rect 12299 5188 12624 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 12728 5148 12756 5179
rect 11379 5120 11744 5148
rect 12360 5120 12756 5148
rect 11379 5117 11391 5120
rect 11333 5111 11391 5117
rect 5813 5083 5871 5089
rect 5813 5049 5825 5083
rect 5859 5049 5871 5083
rect 5813 5043 5871 5049
rect 12360 5024 12388 5120
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 4062 5012 4068 5024
rect 3651 4984 4068 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4249 5015 4307 5021
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 4706 5012 4712 5024
rect 4295 4984 4712 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 5166 5021 5172 5024
rect 5150 5015 5172 5021
rect 5150 4981 5162 5015
rect 5150 4975 5172 4981
rect 5166 4972 5172 4975
rect 5224 4972 5230 5024
rect 5626 4972 5632 5024
rect 5684 4972 5690 5024
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6822 5012 6828 5024
rect 6052 4984 6828 5012
rect 6052 4972 6058 4984
rect 6822 4972 6828 4984
rect 6880 4972 6886 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 8536 4984 8861 5012
rect 8536 4972 8542 4984
rect 8849 4981 8861 4984
rect 8895 4981 8907 5015
rect 8849 4975 8907 4981
rect 9033 5015 9091 5021
rect 9033 4981 9045 5015
rect 9079 5012 9091 5015
rect 9674 5012 9680 5024
rect 9079 4984 9680 5012
rect 9079 4981 9091 4984
rect 9033 4975 9091 4981
rect 9674 4972 9680 4984
rect 9732 4972 9738 5024
rect 12342 4972 12348 5024
rect 12400 4972 12406 5024
rect 1104 4922 13340 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 13340 4922
rect 1104 4848 13340 4870
rect 2041 4811 2099 4817
rect 2041 4777 2053 4811
rect 2087 4808 2099 4811
rect 2130 4808 2136 4820
rect 2087 4780 2136 4808
rect 2087 4777 2099 4780
rect 2041 4771 2099 4777
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 2225 4811 2283 4817
rect 2225 4777 2237 4811
rect 2271 4808 2283 4811
rect 3326 4808 3332 4820
rect 2271 4780 3332 4808
rect 2271 4777 2283 4780
rect 2225 4771 2283 4777
rect 3326 4768 3332 4780
rect 3384 4768 3390 4820
rect 3786 4768 3792 4820
rect 3844 4808 3850 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 3844 4780 3893 4808
rect 3844 4768 3850 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 6638 4808 6644 4820
rect 6227 4780 6644 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 6638 4768 6644 4780
rect 6696 4768 6702 4820
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 10100 4780 10916 4808
rect 10100 4768 10106 4780
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 3694 4740 3700 4752
rect 2639 4712 3700 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 3694 4700 3700 4712
rect 3752 4700 3758 4752
rect 4617 4743 4675 4749
rect 4617 4709 4629 4743
rect 4663 4740 4675 4743
rect 4663 4712 5212 4740
rect 4663 4709 4675 4712
rect 4617 4703 4675 4709
rect 5184 4684 5212 4712
rect 6454 4700 6460 4752
rect 6512 4740 6518 4752
rect 6733 4743 6791 4749
rect 6733 4740 6745 4743
rect 6512 4712 6745 4740
rect 6512 4700 6518 4712
rect 6733 4709 6745 4712
rect 6779 4709 6791 4743
rect 10888 4740 10916 4780
rect 10962 4768 10968 4820
rect 11020 4808 11026 4820
rect 12253 4811 12311 4817
rect 12253 4808 12265 4811
rect 11020 4780 12265 4808
rect 11020 4768 11026 4780
rect 12253 4777 12265 4780
rect 12299 4777 12311 4811
rect 12253 4771 12311 4777
rect 11885 4743 11943 4749
rect 11885 4740 11897 4743
rect 10888 4712 11897 4740
rect 6733 4703 6791 4709
rect 11885 4709 11897 4712
rect 11931 4709 11943 4743
rect 11885 4703 11943 4709
rect 4706 4632 4712 4684
rect 4764 4672 4770 4684
rect 4764 4644 5120 4672
rect 4764 4632 4770 4644
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3973 4607 4031 4613
rect 3973 4604 3985 4607
rect 3200 4576 3985 4604
rect 3200 4564 3206 4576
rect 3973 4573 3985 4576
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 4890 4564 4896 4616
rect 4948 4564 4954 4616
rect 5092 4613 5120 4644
rect 5166 4632 5172 4684
rect 5224 4632 5230 4684
rect 6472 4644 6776 4672
rect 6472 4613 6500 4644
rect 6748 4613 6776 4644
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 7892 4644 8524 4672
rect 7892 4632 7898 4644
rect 8496 4613 8524 4644
rect 9674 4632 9680 4684
rect 9732 4632 9738 4684
rect 5077 4607 5135 4613
rect 5077 4573 5089 4607
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 6457 4607 6515 4613
rect 6457 4573 6469 4607
rect 6503 4573 6515 4607
rect 6457 4567 6515 4573
rect 6549 4607 6607 4613
rect 6549 4573 6561 4607
rect 6595 4573 6607 4607
rect 6549 4567 6607 4573
rect 6733 4607 6791 4613
rect 6733 4573 6745 4607
rect 6779 4604 6791 4607
rect 8481 4607 8539 4613
rect 6779 4576 8064 4604
rect 6779 4573 6791 4576
rect 6733 4567 6791 4573
rect 2225 4539 2283 4545
rect 2225 4505 2237 4539
rect 2271 4536 2283 4539
rect 2406 4536 2412 4548
rect 2271 4508 2412 4536
rect 2271 4505 2283 4508
rect 2225 4499 2283 4505
rect 2406 4496 2412 4508
rect 2464 4496 2470 4548
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 4617 4539 4675 4545
rect 4617 4536 4629 4539
rect 4120 4508 4629 4536
rect 4120 4496 4126 4508
rect 4617 4505 4629 4508
rect 4663 4536 4675 4539
rect 5994 4536 6000 4548
rect 4663 4508 6000 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 5994 4496 6000 4508
rect 6052 4496 6058 4548
rect 6178 4496 6184 4548
rect 6236 4496 6242 4548
rect 6564 4536 6592 4567
rect 8036 4548 8064 4576
rect 8481 4573 8493 4607
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4573 8631 4607
rect 8573 4567 8631 4573
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 6472 4508 6592 4536
rect 6472 4480 6500 4508
rect 7834 4496 7840 4548
rect 7892 4496 7898 4548
rect 8018 4496 8024 4548
rect 8076 4536 8082 4548
rect 8588 4536 8616 4567
rect 8076 4508 8616 4536
rect 9416 4536 9444 4567
rect 10778 4564 10784 4616
rect 10836 4564 10842 4616
rect 11238 4564 11244 4616
rect 11296 4604 11302 4616
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 11296 4576 11529 4604
rect 11296 4564 11302 4576
rect 11517 4573 11529 4576
rect 11563 4573 11575 4607
rect 11517 4567 11575 4573
rect 11698 4564 11704 4616
rect 11756 4564 11762 4616
rect 12342 4613 12348 4616
rect 12337 4604 12348 4613
rect 12303 4576 12348 4604
rect 12337 4567 12348 4576
rect 12342 4564 12348 4567
rect 12400 4564 12406 4616
rect 9582 4536 9588 4548
rect 9416 4508 9588 4536
rect 8076 4496 8082 4508
rect 9582 4496 9588 4508
rect 9640 4496 9646 4548
rect 11425 4539 11483 4545
rect 11425 4505 11437 4539
rect 11471 4505 11483 4539
rect 11425 4499 11483 4505
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 5316 4440 5457 4468
rect 5316 4428 5322 4440
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 6365 4471 6423 4477
rect 6365 4437 6377 4471
rect 6411 4468 6423 4471
rect 6454 4468 6460 4480
rect 6411 4440 6460 4468
rect 6411 4437 6423 4440
rect 6365 4431 6423 4437
rect 6454 4428 6460 4440
rect 6512 4428 6518 4480
rect 8110 4428 8116 4480
rect 8168 4468 8174 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 8168 4440 8217 4468
rect 8168 4428 8174 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 8294 4428 8300 4480
rect 8352 4428 8358 4480
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 11440 4468 11468 4499
rect 9364 4440 11468 4468
rect 9364 4428 9370 4440
rect 1104 4378 13340 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 13340 4378
rect 1104 4304 13340 4326
rect 3694 4224 3700 4276
rect 3752 4264 3758 4276
rect 7834 4264 7840 4276
rect 3752 4236 7840 4264
rect 3752 4224 3758 4236
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 7926 4224 7932 4276
rect 7984 4264 7990 4276
rect 8113 4267 8171 4273
rect 8113 4264 8125 4267
rect 7984 4236 8125 4264
rect 7984 4224 7990 4236
rect 8113 4233 8125 4236
rect 8159 4233 8171 4267
rect 9030 4264 9036 4276
rect 8113 4227 8171 4233
rect 8588 4236 9036 4264
rect 5718 4196 5724 4208
rect 4724 4168 5724 4196
rect 4724 4137 4752 4168
rect 5718 4156 5724 4168
rect 5776 4156 5782 4208
rect 8588 4205 8616 4236
rect 9030 4224 9036 4236
rect 9088 4224 9094 4276
rect 8573 4199 8631 4205
rect 8573 4165 8585 4199
rect 8619 4165 8631 4199
rect 8573 4159 8631 4165
rect 8789 4199 8847 4205
rect 8789 4165 8801 4199
rect 8835 4196 8847 4199
rect 8835 4168 10364 4196
rect 8835 4165 8847 4168
rect 8789 4159 8847 4165
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4097 4767 4131
rect 4709 4091 4767 4097
rect 5491 4131 5549 4137
rect 5491 4097 5503 4131
rect 5537 4128 5549 4131
rect 5626 4128 5632 4140
rect 5537 4100 5632 4128
rect 5537 4097 5549 4100
rect 5491 4091 5549 4097
rect 5626 4088 5632 4100
rect 5684 4088 5690 4140
rect 5810 4088 5816 4140
rect 5868 4128 5874 4140
rect 5997 4131 6055 4137
rect 5997 4128 6009 4131
rect 5868 4100 6009 4128
rect 5868 4088 5874 4100
rect 5997 4097 6009 4100
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6178 4088 6184 4140
rect 6236 4128 6242 4140
rect 6822 4128 6828 4140
rect 6236 4100 6828 4128
rect 6236 4088 6242 4100
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 9217 4131 9275 4137
rect 9217 4128 9229 4131
rect 6932 4100 9229 4128
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 3881 4063 3939 4069
rect 3881 4060 3893 4063
rect 2832 4032 3893 4060
rect 2832 4020 2838 4032
rect 3881 4029 3893 4032
rect 3927 4060 3939 4063
rect 4433 4063 4491 4069
rect 3927 4032 4384 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 4356 3924 4384 4032
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 4798 4060 4804 4072
rect 4479 4032 4804 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 4893 4063 4951 4069
rect 4893 4029 4905 4063
rect 4939 4060 4951 4063
rect 4985 4063 5043 4069
rect 4985 4060 4997 4063
rect 4939 4032 4997 4060
rect 4939 4029 4951 4032
rect 4893 4023 4951 4029
rect 4985 4029 4997 4032
rect 5031 4029 5043 4063
rect 4985 4023 5043 4029
rect 5350 4020 5356 4072
rect 5408 4020 5414 4072
rect 6932 4060 6960 4100
rect 9217 4097 9229 4100
rect 9263 4097 9275 4131
rect 9953 4131 10011 4137
rect 9953 4128 9965 4131
rect 9217 4091 9275 4097
rect 9324 4100 9965 4128
rect 5460 4032 6960 4060
rect 5460 3924 5488 4032
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8352 4032 8493 4060
rect 8352 4020 8358 4032
rect 8481 4029 8493 4032
rect 8527 4060 8539 4063
rect 9324 4060 9352 4100
rect 9953 4097 9965 4100
rect 9999 4097 10011 4131
rect 9953 4091 10011 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 10226 4128 10232 4140
rect 10183 4100 10232 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10336 4137 10364 4168
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 8527 4032 9352 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9456 4032 9505 4060
rect 9456 4020 9462 4032
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 10612 4060 10640 4091
rect 10778 4088 10784 4140
rect 10836 4088 10842 4140
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 12342 4128 12348 4140
rect 10919 4100 12348 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 10888 4060 10916 4091
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 9493 4023 9551 4029
rect 9646 4032 10916 4060
rect 5902 3952 5908 4004
rect 5960 3992 5966 4004
rect 6089 3995 6147 4001
rect 6089 3992 6101 3995
rect 5960 3964 6101 3992
rect 5960 3952 5966 3964
rect 6089 3961 6101 3964
rect 6135 3961 6147 3995
rect 6089 3955 6147 3961
rect 8570 3952 8576 4004
rect 8628 3992 8634 4004
rect 9646 3992 9674 4032
rect 8628 3964 9674 3992
rect 8628 3952 8634 3964
rect 4356 3896 5488 3924
rect 5534 3884 5540 3936
rect 5592 3884 5598 3936
rect 7926 3884 7932 3936
rect 7984 3884 7990 3936
rect 8110 3884 8116 3936
rect 8168 3884 8174 3936
rect 8754 3884 8760 3936
rect 8812 3884 8818 3936
rect 8938 3884 8944 3936
rect 8996 3884 9002 3936
rect 10502 3884 10508 3936
rect 10560 3884 10566 3936
rect 1104 3834 13340 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 13340 3834
rect 1104 3760 13340 3782
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 4856 3692 5089 3720
rect 4856 3680 4862 3692
rect 5077 3689 5089 3692
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 5350 3680 5356 3732
rect 5408 3720 5414 3732
rect 5813 3723 5871 3729
rect 5813 3720 5825 3723
rect 5408 3692 5825 3720
rect 5408 3680 5414 3692
rect 5813 3689 5825 3692
rect 5859 3689 5871 3723
rect 5813 3683 5871 3689
rect 6454 3680 6460 3732
rect 6512 3680 6518 3732
rect 8297 3723 8355 3729
rect 8297 3689 8309 3723
rect 8343 3720 8355 3723
rect 8754 3720 8760 3732
rect 8343 3692 8760 3720
rect 8343 3689 8355 3692
rect 8297 3683 8355 3689
rect 8754 3680 8760 3692
rect 8812 3680 8818 3732
rect 8938 3680 8944 3732
rect 8996 3720 9002 3732
rect 9198 3723 9256 3729
rect 9198 3720 9210 3723
rect 8996 3692 9210 3720
rect 8996 3680 9002 3692
rect 9198 3689 9210 3692
rect 9244 3689 9256 3723
rect 9198 3683 9256 3689
rect 10226 3680 10232 3732
rect 10284 3720 10290 3732
rect 10689 3723 10747 3729
rect 10689 3720 10701 3723
rect 10284 3692 10701 3720
rect 10284 3680 10290 3692
rect 10689 3689 10701 3692
rect 10735 3689 10747 3723
rect 10689 3683 10747 3689
rect 12618 3680 12624 3732
rect 12676 3720 12682 3732
rect 12805 3723 12863 3729
rect 12805 3720 12817 3723
rect 12676 3692 12817 3720
rect 12676 3680 12682 3692
rect 12805 3689 12817 3692
rect 12851 3689 12863 3723
rect 12805 3683 12863 3689
rect 4614 3612 4620 3664
rect 4672 3612 4678 3664
rect 4985 3655 5043 3661
rect 4985 3621 4997 3655
rect 5031 3652 5043 3655
rect 5031 3624 6040 3652
rect 5031 3621 5043 3624
rect 4985 3615 5043 3621
rect 4632 3584 4660 3612
rect 6012 3596 6040 3624
rect 4709 3587 4767 3593
rect 4709 3584 4721 3587
rect 4632 3556 4721 3584
rect 4709 3553 4721 3556
rect 4755 3553 4767 3587
rect 4709 3547 4767 3553
rect 5258 3544 5264 3596
rect 5316 3544 5322 3596
rect 5445 3587 5503 3593
rect 5445 3553 5457 3587
rect 5491 3584 5503 3587
rect 5902 3584 5908 3596
rect 5491 3556 5908 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 5994 3544 6000 3596
rect 6052 3544 6058 3596
rect 8018 3584 8024 3596
rect 6104 3556 8024 3584
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4798 3516 4804 3528
rect 4663 3488 4804 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4798 3476 4804 3488
rect 4856 3476 4862 3528
rect 5350 3476 5356 3528
rect 5408 3476 5414 3528
rect 5534 3476 5540 3528
rect 5592 3476 5598 3528
rect 6104 3525 6132 3556
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8938 3544 8944 3596
rect 8996 3584 9002 3596
rect 9582 3584 9588 3596
rect 8996 3556 9588 3584
rect 8996 3544 9002 3556
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 6178 3516 6184 3528
rect 6135 3488 6184 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 6638 3476 6644 3528
rect 6696 3476 6702 3528
rect 6822 3476 6828 3528
rect 6880 3476 6886 3528
rect 6914 3476 6920 3528
rect 6972 3476 6978 3528
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7190 3516 7196 3528
rect 7147 3488 7196 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7190 3476 7196 3488
rect 7248 3476 7254 3528
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 5552 3448 5580 3476
rect 6733 3451 6791 3457
rect 6733 3448 6745 3451
rect 5552 3420 6745 3448
rect 6733 3417 6745 3420
rect 6779 3417 6791 3451
rect 6840 3448 6868 3476
rect 8220 3448 8248 3479
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8389 3519 8447 3525
rect 8389 3516 8401 3519
rect 8352 3488 8401 3516
rect 8352 3476 8358 3488
rect 8389 3485 8401 3488
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 12986 3476 12992 3528
rect 13044 3476 13050 3528
rect 10502 3448 10508 3460
rect 6840 3420 8800 3448
rect 10442 3420 10508 3448
rect 6733 3411 6791 3417
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 6638 3380 6644 3392
rect 5868 3352 6644 3380
rect 5868 3340 5874 3352
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 7006 3340 7012 3392
rect 7064 3340 7070 3392
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 8665 3383 8723 3389
rect 8665 3380 8677 3383
rect 8628 3352 8677 3380
rect 8628 3340 8634 3352
rect 8665 3349 8677 3352
rect 8711 3349 8723 3383
rect 8772 3380 8800 3420
rect 10502 3408 10508 3420
rect 10560 3408 10566 3460
rect 10226 3380 10232 3392
rect 8772 3352 10232 3380
rect 8665 3343 8723 3349
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 1104 3290 13340 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 13340 3290
rect 1104 3216 13340 3238
rect 5350 3136 5356 3188
rect 5408 3176 5414 3188
rect 6089 3179 6147 3185
rect 6089 3176 6101 3179
rect 5408 3148 6101 3176
rect 5408 3136 5414 3148
rect 6089 3145 6101 3148
rect 6135 3145 6147 3179
rect 6089 3139 6147 3145
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 8113 3179 8171 3185
rect 8113 3176 8125 3179
rect 8076 3148 8125 3176
rect 8076 3136 8082 3148
rect 8113 3145 8125 3148
rect 8159 3145 8171 3179
rect 8113 3139 8171 3145
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 6914 3108 6920 3120
rect 4672 3080 6920 3108
rect 4672 3068 4678 3080
rect 6914 3068 6920 3080
rect 6972 3068 6978 3120
rect 8570 3068 8576 3120
rect 8628 3068 8634 3120
rect 9582 3068 9588 3120
rect 9640 3108 9646 3120
rect 9640 3080 9904 3108
rect 9640 3068 9646 3080
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3009 5595 3043
rect 5537 3003 5595 3009
rect 5552 2904 5580 3003
rect 5994 3000 6000 3052
rect 6052 3000 6058 3052
rect 6178 3000 6184 3052
rect 6236 3000 6242 3052
rect 6454 3000 6460 3052
rect 6512 3040 6518 3052
rect 6733 3043 6791 3049
rect 6733 3040 6745 3043
rect 6512 3012 6745 3040
rect 6512 3000 6518 3012
rect 6733 3009 6745 3012
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 9876 3049 9904 3080
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7616 3012 7849 3040
rect 7616 3000 7622 3012
rect 7837 3009 7849 3012
rect 7883 3009 7895 3043
rect 7837 3003 7895 3009
rect 9861 3043 9919 3049
rect 9861 3009 9873 3043
rect 9907 3009 9919 3043
rect 9861 3003 9919 3009
rect 5629 2975 5687 2981
rect 5629 2941 5641 2975
rect 5675 2972 5687 2975
rect 7006 2972 7012 2984
rect 5675 2944 7012 2972
rect 5675 2941 5687 2944
rect 5629 2935 5687 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 7926 2932 7932 2984
rect 7984 2972 7990 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 7984 2944 9597 2972
rect 7984 2932 7990 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 6546 2904 6552 2916
rect 5552 2876 6552 2904
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 5810 2796 5816 2848
rect 5868 2796 5874 2848
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7285 2839 7343 2845
rect 7285 2836 7297 2839
rect 7156 2808 7297 2836
rect 7156 2796 7162 2808
rect 7285 2805 7297 2808
rect 7331 2805 7343 2839
rect 7285 2799 7343 2805
rect 7742 2796 7748 2848
rect 7800 2796 7806 2848
rect 1104 2746 13340 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 13340 2746
rect 1104 2672 13340 2694
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 5442 2632 5448 2644
rect 5123 2604 5448 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 7190 2632 7196 2644
rect 5736 2604 7196 2632
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 5736 2496 5764 2604
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 7524 2604 8217 2632
rect 7524 2592 7530 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 4856 2468 5764 2496
rect 4856 2456 4862 2468
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 5736 2428 5764 2468
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 6181 2499 6239 2505
rect 6181 2496 6193 2499
rect 5868 2468 6193 2496
rect 5868 2456 5874 2468
rect 6181 2465 6193 2468
rect 6227 2465 6239 2499
rect 6181 2459 6239 2465
rect 6457 2499 6515 2505
rect 6457 2465 6469 2499
rect 6503 2496 6515 2499
rect 8938 2496 8944 2508
rect 6503 2468 8944 2496
rect 6503 2465 6515 2468
rect 6457 2459 6515 2465
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5736 2400 5917 2428
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 6730 2320 6736 2372
rect 6788 2320 6794 2372
rect 7742 2320 7748 2372
rect 7800 2320 7806 2372
rect 1104 2202 13340 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 13340 2202
rect 1104 2128 13340 2150
<< via1 >>
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 8392 13948 8444 14000
rect 5264 13923 5316 13932
rect 5264 13889 5273 13923
rect 5273 13889 5307 13923
rect 5307 13889 5316 13923
rect 5264 13880 5316 13889
rect 5816 13880 5868 13932
rect 6460 13880 6512 13932
rect 7104 13880 7156 13932
rect 7748 13880 7800 13932
rect 9128 13880 9180 13932
rect 9680 13880 9732 13932
rect 8300 13812 8352 13864
rect 9404 13812 9456 13864
rect 4712 13744 4764 13796
rect 6644 13744 6696 13796
rect 9772 13744 9824 13796
rect 9864 13744 9916 13796
rect 5908 13719 5960 13728
rect 5908 13685 5917 13719
rect 5917 13685 5951 13719
rect 5951 13685 5960 13719
rect 5908 13676 5960 13685
rect 6736 13719 6788 13728
rect 6736 13685 6745 13719
rect 6745 13685 6779 13719
rect 6779 13685 6788 13719
rect 6736 13676 6788 13685
rect 7196 13676 7248 13728
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 5816 13472 5868 13524
rect 6736 13472 6788 13524
rect 3608 13404 3660 13456
rect 6460 13404 6512 13456
rect 4804 13336 4856 13388
rect 5264 13336 5316 13388
rect 5908 13336 5960 13388
rect 7012 13336 7064 13388
rect 8300 13472 8352 13524
rect 9864 13404 9916 13456
rect 3056 13200 3108 13252
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 5632 13268 5684 13320
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 6644 13311 6696 13320
rect 6644 13277 6653 13311
rect 6653 13277 6687 13311
rect 6687 13277 6696 13311
rect 6644 13268 6696 13277
rect 9956 13336 10008 13388
rect 7196 13268 7248 13320
rect 8208 13268 8260 13320
rect 3792 13132 3844 13184
rect 5724 13200 5776 13252
rect 4252 13132 4304 13184
rect 6276 13175 6328 13184
rect 6276 13141 6285 13175
rect 6285 13141 6319 13175
rect 6319 13141 6328 13175
rect 6276 13132 6328 13141
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 8116 13243 8168 13252
rect 8116 13209 8125 13243
rect 8125 13209 8159 13243
rect 8159 13209 8168 13243
rect 8116 13200 8168 13209
rect 9496 13268 9548 13320
rect 10048 13200 10100 13252
rect 7840 13132 7892 13184
rect 9680 13132 9732 13184
rect 10416 13132 10468 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 4988 12928 5040 12980
rect 6920 12928 6972 12980
rect 7196 12971 7248 12980
rect 7196 12937 7205 12971
rect 7205 12937 7239 12971
rect 7239 12937 7248 12971
rect 7196 12928 7248 12937
rect 3792 12835 3844 12844
rect 3792 12801 3801 12835
rect 3801 12801 3835 12835
rect 3835 12801 3844 12835
rect 3792 12792 3844 12801
rect 4252 12835 4304 12844
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 4528 12724 4580 12776
rect 4712 12835 4764 12844
rect 4712 12801 4721 12835
rect 4721 12801 4755 12835
rect 4755 12801 4764 12835
rect 4712 12792 4764 12801
rect 4344 12699 4396 12708
rect 4344 12665 4353 12699
rect 4353 12665 4387 12699
rect 4387 12665 4396 12699
rect 4344 12656 4396 12665
rect 4712 12656 4764 12708
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 5264 12792 5316 12844
rect 5632 12792 5684 12844
rect 6552 12792 6604 12844
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7656 12835 7708 12844
rect 7656 12801 7665 12835
rect 7665 12801 7699 12835
rect 7699 12801 7708 12835
rect 7656 12792 7708 12801
rect 7748 12835 7800 12844
rect 7748 12801 7757 12835
rect 7757 12801 7791 12835
rect 7791 12801 7800 12835
rect 7748 12792 7800 12801
rect 9680 12928 9732 12980
rect 9956 12971 10008 12980
rect 9956 12937 9965 12971
rect 9965 12937 9999 12971
rect 9999 12937 10008 12971
rect 9956 12928 10008 12937
rect 7472 12724 7524 12776
rect 6368 12656 6420 12708
rect 7380 12699 7432 12708
rect 7380 12665 7389 12699
rect 7389 12665 7423 12699
rect 7423 12665 7432 12699
rect 7380 12656 7432 12665
rect 3516 12631 3568 12640
rect 3516 12597 3525 12631
rect 3525 12597 3559 12631
rect 3559 12597 3568 12631
rect 3516 12588 3568 12597
rect 5080 12588 5132 12640
rect 5172 12631 5224 12640
rect 5172 12597 5181 12631
rect 5181 12597 5215 12631
rect 5215 12597 5224 12631
rect 5172 12588 5224 12597
rect 6736 12631 6788 12640
rect 6736 12597 6745 12631
rect 6745 12597 6779 12631
rect 6779 12597 6788 12631
rect 6736 12588 6788 12597
rect 6920 12588 6972 12640
rect 8852 12792 8904 12844
rect 9496 12860 9548 12912
rect 8300 12724 8352 12776
rect 8392 12656 8444 12708
rect 9404 12835 9456 12844
rect 9404 12801 9413 12835
rect 9413 12801 9447 12835
rect 9447 12801 9456 12835
rect 9404 12792 9456 12801
rect 9864 12835 9916 12844
rect 9864 12801 9873 12835
rect 9873 12801 9907 12835
rect 9907 12801 9916 12835
rect 9864 12792 9916 12801
rect 10048 12835 10100 12844
rect 10048 12801 10057 12835
rect 10057 12801 10091 12835
rect 10091 12801 10100 12835
rect 10048 12792 10100 12801
rect 11244 12792 11296 12844
rect 9220 12631 9272 12640
rect 9220 12597 9229 12631
rect 9229 12597 9263 12631
rect 9263 12597 9272 12631
rect 9220 12588 9272 12597
rect 9496 12631 9548 12640
rect 9496 12597 9505 12631
rect 9505 12597 9539 12631
rect 9539 12597 9548 12631
rect 9496 12588 9548 12597
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 3056 12427 3108 12436
rect 3056 12393 3065 12427
rect 3065 12393 3099 12427
rect 3099 12393 3108 12427
rect 3056 12384 3108 12393
rect 3608 12384 3660 12436
rect 4068 12427 4120 12436
rect 4068 12393 4077 12427
rect 4077 12393 4111 12427
rect 4111 12393 4120 12427
rect 4068 12384 4120 12393
rect 6276 12384 6328 12436
rect 7012 12384 7064 12436
rect 11336 12427 11388 12436
rect 11336 12393 11345 12427
rect 11345 12393 11379 12427
rect 11379 12393 11388 12427
rect 11336 12384 11388 12393
rect 3792 12248 3844 12300
rect 4344 12248 4396 12300
rect 4528 12291 4580 12300
rect 4528 12257 4537 12291
rect 4537 12257 4571 12291
rect 4571 12257 4580 12291
rect 4528 12248 4580 12257
rect 4252 12223 4304 12232
rect 4252 12189 4261 12223
rect 4261 12189 4295 12223
rect 4295 12189 4304 12223
rect 4252 12180 4304 12189
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 5080 12248 5132 12300
rect 5908 12248 5960 12300
rect 3516 12112 3568 12164
rect 4160 12112 4212 12164
rect 8300 12359 8352 12368
rect 8300 12325 8309 12359
rect 8309 12325 8343 12359
rect 8343 12325 8352 12359
rect 8300 12316 8352 12325
rect 9128 12316 9180 12368
rect 7840 12291 7892 12300
rect 7840 12257 7849 12291
rect 7849 12257 7883 12291
rect 7883 12257 7892 12291
rect 7840 12248 7892 12257
rect 6828 12180 6880 12232
rect 7472 12180 7524 12232
rect 8484 12248 8536 12300
rect 8116 12180 8168 12232
rect 8576 12180 8628 12232
rect 9128 12223 9180 12232
rect 9128 12189 9137 12223
rect 9137 12189 9171 12223
rect 9171 12189 9180 12223
rect 9128 12180 9180 12189
rect 9220 12223 9272 12232
rect 9220 12189 9229 12223
rect 9229 12189 9263 12223
rect 9263 12189 9272 12223
rect 9220 12180 9272 12189
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 9864 12180 9916 12232
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 10416 12223 10468 12232
rect 10416 12189 10425 12223
rect 10425 12189 10459 12223
rect 10459 12189 10468 12223
rect 10416 12180 10468 12189
rect 10600 12180 10652 12232
rect 3332 12044 3384 12096
rect 4436 12044 4488 12096
rect 5356 12044 5408 12096
rect 5908 12044 5960 12096
rect 7932 12044 7984 12096
rect 9036 12044 9088 12096
rect 9128 12044 9180 12096
rect 9956 12112 10008 12164
rect 10140 12112 10192 12164
rect 9496 12044 9548 12096
rect 10048 12044 10100 12096
rect 10876 12180 10928 12232
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11796 12223 11848 12232
rect 11796 12189 11805 12223
rect 11805 12189 11839 12223
rect 11839 12189 11848 12223
rect 11796 12180 11848 12189
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 4252 11840 4304 11892
rect 4344 11840 4396 11892
rect 4896 11840 4948 11892
rect 3516 11772 3568 11824
rect 4988 11772 5040 11824
rect 5724 11840 5776 11892
rect 11796 11840 11848 11892
rect 12624 11840 12676 11892
rect 3792 11704 3844 11756
rect 4068 11747 4120 11756
rect 4068 11713 4077 11747
rect 4077 11713 4111 11747
rect 4111 11713 4120 11747
rect 4068 11704 4120 11713
rect 4160 11747 4212 11756
rect 4160 11713 4169 11747
rect 4169 11713 4203 11747
rect 4203 11713 4212 11747
rect 4160 11704 4212 11713
rect 4804 11704 4856 11756
rect 5080 11747 5132 11756
rect 5080 11713 5089 11747
rect 5089 11713 5123 11747
rect 5123 11713 5132 11747
rect 5080 11704 5132 11713
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 5264 11747 5316 11756
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 5908 11772 5960 11824
rect 5632 11704 5684 11756
rect 6184 11704 6236 11756
rect 6644 11704 6696 11756
rect 7932 11747 7984 11756
rect 7932 11713 7941 11747
rect 7941 11713 7975 11747
rect 7975 11713 7984 11747
rect 7932 11704 7984 11713
rect 8484 11772 8536 11824
rect 12532 11815 12584 11824
rect 12532 11781 12541 11815
rect 12541 11781 12575 11815
rect 12575 11781 12584 11815
rect 12532 11772 12584 11781
rect 8852 11704 8904 11756
rect 9128 11704 9180 11756
rect 6460 11636 6512 11688
rect 8392 11636 8444 11688
rect 8576 11636 8628 11688
rect 9312 11747 9364 11756
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 9680 11704 9732 11756
rect 11060 11704 11112 11756
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 10876 11636 10928 11688
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 4712 11568 4764 11620
rect 5172 11568 5224 11620
rect 6368 11568 6420 11620
rect 4620 11500 4672 11552
rect 5356 11500 5408 11552
rect 5632 11543 5684 11552
rect 5632 11509 5641 11543
rect 5641 11509 5675 11543
rect 5675 11509 5684 11543
rect 5632 11500 5684 11509
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 8484 11500 8536 11509
rect 8944 11500 8996 11552
rect 12256 11500 12308 11552
rect 12716 11500 12768 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 4068 11296 4120 11348
rect 4712 11296 4764 11348
rect 4896 11296 4948 11348
rect 5172 11228 5224 11280
rect 5080 11160 5132 11212
rect 3516 10956 3568 11008
rect 3976 11024 4028 11076
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5632 11160 5684 11212
rect 11060 11296 11112 11348
rect 7932 11160 7984 11212
rect 11244 11160 11296 11212
rect 4712 11067 4764 11076
rect 4712 11033 4721 11067
rect 4721 11033 4755 11067
rect 4755 11033 4764 11067
rect 4712 11024 4764 11033
rect 8392 11092 8444 11144
rect 9496 11092 9548 11144
rect 9680 11092 9732 11144
rect 10876 11092 10928 11144
rect 12716 11160 12768 11212
rect 12808 11092 12860 11144
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 6276 11024 6328 11076
rect 12440 11067 12492 11076
rect 12440 11033 12449 11067
rect 12449 11033 12483 11067
rect 12483 11033 12492 11067
rect 12440 11024 12492 11033
rect 5264 10956 5316 11008
rect 5448 10999 5500 11008
rect 5448 10965 5457 10999
rect 5457 10965 5491 10999
rect 5491 10965 5500 10999
rect 5448 10956 5500 10965
rect 5908 10999 5960 11008
rect 5908 10965 5917 10999
rect 5917 10965 5951 10999
rect 5951 10965 5960 10999
rect 5908 10956 5960 10965
rect 8024 10956 8076 11008
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 10324 10956 10376 11008
rect 11980 10999 12032 11008
rect 11980 10965 11989 10999
rect 11989 10965 12023 10999
rect 12023 10965 12032 10999
rect 11980 10956 12032 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 11888 10752 11940 10804
rect 3884 10684 3936 10736
rect 5908 10684 5960 10736
rect 5264 10616 5316 10668
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 5724 10616 5776 10668
rect 1676 10548 1728 10600
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 2780 10412 2832 10464
rect 5816 10548 5868 10600
rect 8484 10684 8536 10736
rect 9220 10684 9272 10736
rect 11244 10684 11296 10736
rect 11980 10684 12032 10736
rect 12624 10684 12676 10736
rect 6552 10616 6604 10668
rect 7472 10616 7524 10668
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 7380 10548 7432 10600
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9496 10616 9548 10668
rect 9680 10659 9732 10668
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 12532 10659 12584 10668
rect 8852 10591 8904 10600
rect 8852 10557 8861 10591
rect 8861 10557 8895 10591
rect 8895 10557 8904 10591
rect 8852 10548 8904 10557
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 10324 10591 10376 10600
rect 10324 10557 10333 10591
rect 10333 10557 10367 10591
rect 10367 10557 10376 10591
rect 10324 10548 10376 10557
rect 10232 10480 10284 10532
rect 12532 10625 12541 10659
rect 12541 10625 12575 10659
rect 12575 10625 12584 10659
rect 12532 10616 12584 10625
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 12808 10659 12860 10668
rect 12808 10625 12817 10659
rect 12817 10625 12851 10659
rect 12851 10625 12860 10659
rect 12808 10616 12860 10625
rect 12440 10548 12492 10600
rect 12532 10480 12584 10532
rect 6644 10412 6696 10464
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 7288 10412 7340 10464
rect 8116 10412 8168 10464
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 9864 10455 9916 10464
rect 9864 10421 9873 10455
rect 9873 10421 9907 10455
rect 9907 10421 9916 10455
rect 9864 10412 9916 10421
rect 10692 10412 10744 10464
rect 12624 10412 12676 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3516 10251 3568 10260
rect 3516 10217 3525 10251
rect 3525 10217 3559 10251
rect 3559 10217 3568 10251
rect 3516 10208 3568 10217
rect 3884 10251 3936 10260
rect 3884 10217 3893 10251
rect 3893 10217 3927 10251
rect 3927 10217 3936 10251
rect 3884 10208 3936 10217
rect 4712 10208 4764 10260
rect 6644 10208 6696 10260
rect 2780 10072 2832 10124
rect 3056 10072 3108 10124
rect 3792 10072 3844 10124
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 1676 10047 1728 10056
rect 1676 10013 1685 10047
rect 1685 10013 1719 10047
rect 1719 10013 1728 10047
rect 1676 10004 1728 10013
rect 4068 10004 4120 10056
rect 2044 9979 2096 9988
rect 2044 9945 2053 9979
rect 2053 9945 2087 9979
rect 2087 9945 2096 9979
rect 2044 9936 2096 9945
rect 4712 10004 4764 10056
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 5448 10004 5500 10056
rect 5540 10004 5592 10056
rect 5724 10047 5776 10056
rect 5724 10013 5733 10047
rect 5733 10013 5767 10047
rect 5767 10013 5776 10047
rect 5724 10004 5776 10013
rect 4620 9936 4672 9988
rect 5908 9936 5960 9988
rect 3332 9868 3384 9920
rect 4160 9868 4212 9920
rect 5540 9868 5592 9920
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 6736 10004 6788 10056
rect 8760 10140 8812 10192
rect 8024 10072 8076 10124
rect 7288 10047 7340 10056
rect 7288 10013 7297 10047
rect 7297 10013 7331 10047
rect 7331 10013 7340 10047
rect 7288 10004 7340 10013
rect 7748 10004 7800 10056
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8944 10004 8996 10056
rect 12440 10251 12492 10260
rect 9588 10140 9640 10192
rect 12440 10217 12449 10251
rect 12449 10217 12483 10251
rect 12483 10217 12492 10251
rect 12440 10208 12492 10217
rect 12716 10208 12768 10260
rect 9680 10047 9732 10056
rect 9680 10013 9689 10047
rect 9689 10013 9723 10047
rect 9723 10013 9732 10047
rect 9680 10004 9732 10013
rect 9772 10047 9824 10056
rect 9772 10013 9782 10047
rect 9782 10013 9816 10047
rect 9816 10013 9824 10047
rect 9772 10004 9824 10013
rect 10600 10047 10652 10056
rect 10600 10013 10609 10047
rect 10609 10013 10643 10047
rect 10643 10013 10652 10047
rect 10600 10004 10652 10013
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 10968 10047 11020 10056
rect 7104 9936 7156 9988
rect 9036 9936 9088 9988
rect 9220 9936 9272 9988
rect 10968 10013 10977 10047
rect 10977 10013 11011 10047
rect 11011 10013 11020 10047
rect 10968 10004 11020 10013
rect 11244 10004 11296 10056
rect 12072 10140 12124 10192
rect 12532 10115 12584 10124
rect 12532 10081 12541 10115
rect 12541 10081 12575 10115
rect 12575 10081 12584 10115
rect 12532 10072 12584 10081
rect 12164 10047 12216 10056
rect 12164 10013 12209 10047
rect 12209 10013 12216 10047
rect 12164 10004 12216 10013
rect 12348 10047 12400 10056
rect 12348 10013 12357 10047
rect 12357 10013 12391 10047
rect 12391 10013 12400 10047
rect 12348 10004 12400 10013
rect 12624 10004 12676 10056
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7196 9911 7248 9920
rect 7196 9877 7205 9911
rect 7205 9877 7239 9911
rect 7239 9877 7248 9911
rect 7196 9868 7248 9877
rect 7288 9868 7340 9920
rect 7472 9868 7524 9920
rect 11980 9979 12032 9988
rect 11980 9945 11989 9979
rect 11989 9945 12023 9979
rect 12023 9945 12032 9979
rect 11980 9936 12032 9945
rect 12072 9979 12124 9988
rect 12072 9945 12081 9979
rect 12081 9945 12115 9979
rect 12115 9945 12124 9979
rect 12072 9936 12124 9945
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 1492 9596 1544 9648
rect 1676 9596 1728 9648
rect 2964 9664 3016 9716
rect 3240 9664 3292 9716
rect 4804 9664 4856 9716
rect 2320 9596 2372 9648
rect 4068 9596 4120 9648
rect 4160 9639 4212 9648
rect 4160 9605 4169 9639
rect 4169 9605 4203 9639
rect 4203 9605 4212 9639
rect 4160 9596 4212 9605
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 3884 9528 3936 9580
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 4620 9571 4672 9580
rect 4620 9537 4629 9571
rect 4629 9537 4663 9571
rect 4663 9537 4672 9571
rect 4620 9528 4672 9537
rect 4804 9528 4856 9580
rect 5908 9639 5960 9648
rect 5908 9605 5917 9639
rect 5917 9605 5951 9639
rect 5951 9605 5960 9639
rect 5908 9596 5960 9605
rect 7104 9664 7156 9716
rect 7196 9707 7248 9716
rect 7196 9673 7205 9707
rect 7205 9673 7239 9707
rect 7239 9673 7248 9707
rect 7196 9664 7248 9673
rect 8852 9664 8904 9716
rect 9680 9664 9732 9716
rect 12072 9707 12124 9716
rect 12072 9673 12081 9707
rect 12081 9673 12115 9707
rect 12115 9673 12124 9707
rect 12072 9664 12124 9673
rect 5540 9571 5592 9580
rect 5540 9537 5549 9571
rect 5549 9537 5583 9571
rect 5583 9537 5592 9571
rect 5540 9528 5592 9537
rect 6092 9571 6144 9580
rect 6092 9537 6101 9571
rect 6101 9537 6135 9571
rect 6135 9537 6144 9571
rect 6092 9528 6144 9537
rect 6920 9596 6972 9648
rect 10232 9639 10284 9648
rect 10232 9605 10241 9639
rect 10241 9605 10275 9639
rect 10275 9605 10284 9639
rect 10232 9596 10284 9605
rect 10600 9596 10652 9648
rect 12532 9664 12584 9716
rect 2596 9503 2648 9512
rect 2596 9469 2605 9503
rect 2605 9469 2639 9503
rect 2639 9469 2648 9503
rect 2596 9460 2648 9469
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 5448 9460 5500 9512
rect 6644 9460 6696 9512
rect 2504 9392 2556 9444
rect 2872 9392 2924 9444
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 7288 9528 7340 9580
rect 7380 9571 7432 9580
rect 7380 9537 7389 9571
rect 7389 9537 7423 9571
rect 7423 9537 7432 9571
rect 7380 9528 7432 9537
rect 9312 9571 9364 9580
rect 9312 9537 9321 9571
rect 9321 9537 9355 9571
rect 9355 9537 9364 9571
rect 9312 9528 9364 9537
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 11244 9528 11296 9580
rect 12440 9571 12492 9586
rect 12440 9537 12449 9571
rect 12449 9537 12483 9571
rect 12483 9537 12492 9571
rect 12440 9534 12492 9537
rect 12072 9460 12124 9512
rect 8760 9435 8812 9444
rect 8760 9401 8769 9435
rect 8769 9401 8803 9435
rect 8803 9401 8812 9435
rect 8760 9392 8812 9401
rect 9220 9392 9272 9444
rect 10324 9392 10376 9444
rect 12164 9392 12216 9444
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 12624 9460 12676 9512
rect 12808 9392 12860 9444
rect 3056 9324 3108 9376
rect 3332 9324 3384 9376
rect 4528 9324 4580 9376
rect 4712 9324 4764 9376
rect 6276 9324 6328 9376
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 9772 9324 9824 9376
rect 10968 9324 11020 9376
rect 12716 9324 12768 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2504 8984 2556 9036
rect 2964 9052 3016 9104
rect 6092 9120 6144 9172
rect 6828 9120 6880 9172
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 10968 9120 11020 9172
rect 12624 9120 12676 9172
rect 12808 9163 12860 9172
rect 12808 9129 12817 9163
rect 12817 9129 12851 9163
rect 12851 9129 12860 9163
rect 12808 9120 12860 9129
rect 7196 9052 7248 9104
rect 2596 8916 2648 8968
rect 2872 9027 2924 9036
rect 2872 8993 2881 9027
rect 2881 8993 2915 9027
rect 2915 8993 2924 9027
rect 2872 8984 2924 8993
rect 3608 8916 3660 8968
rect 4620 8916 4672 8968
rect 4712 8916 4764 8968
rect 5448 8916 5500 8968
rect 6276 8959 6328 8968
rect 6276 8925 6285 8959
rect 6285 8925 6319 8959
rect 6319 8925 6328 8959
rect 6276 8916 6328 8925
rect 8392 8984 8444 9036
rect 6644 8959 6696 8968
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 9220 8959 9272 8968
rect 9220 8925 9229 8959
rect 9229 8925 9263 8959
rect 9263 8925 9272 8959
rect 9220 8916 9272 8925
rect 9864 8916 9916 8968
rect 11980 8916 12032 8968
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 5264 8848 5316 8900
rect 2228 8780 2280 8832
rect 2596 8780 2648 8832
rect 4712 8780 4764 8832
rect 6736 8780 6788 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2320 8576 2372 8628
rect 2412 8508 2464 8560
rect 2872 8508 2924 8560
rect 3608 8619 3660 8628
rect 3608 8585 3617 8619
rect 3617 8585 3651 8619
rect 3651 8585 3660 8619
rect 3608 8576 3660 8585
rect 4252 8576 4304 8628
rect 4988 8576 5040 8628
rect 5540 8440 5592 8492
rect 6552 8508 6604 8560
rect 10324 8440 10376 8492
rect 12624 8483 12676 8492
rect 12624 8449 12633 8483
rect 12633 8449 12667 8483
rect 12667 8449 12676 8483
rect 12624 8440 12676 8449
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 1860 8415 1912 8424
rect 1860 8381 1869 8415
rect 1869 8381 1903 8415
rect 1903 8381 1912 8415
rect 1860 8372 1912 8381
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 4620 8372 4672 8424
rect 4896 8372 4948 8424
rect 5448 8372 5500 8424
rect 10968 8372 11020 8424
rect 11060 8372 11112 8424
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 3148 8236 3200 8288
rect 5540 8236 5592 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 2228 8075 2280 8084
rect 2228 8041 2237 8075
rect 2237 8041 2271 8075
rect 2271 8041 2280 8075
rect 2228 8032 2280 8041
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 2872 8032 2924 8084
rect 4988 8032 5040 8084
rect 5356 8032 5408 8084
rect 6000 8032 6052 8084
rect 7748 8032 7800 8084
rect 10416 8032 10468 8084
rect 12072 8032 12124 8084
rect 1860 7964 1912 8016
rect 2780 7964 2832 8016
rect 1584 7828 1636 7880
rect 2596 7828 2648 7880
rect 3148 7828 3200 7880
rect 3976 7964 4028 8016
rect 6276 7896 6328 7948
rect 9404 7896 9456 7948
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8944 7828 8996 7880
rect 12716 7871 12768 7880
rect 12716 7837 12725 7871
rect 12725 7837 12759 7871
rect 12759 7837 12768 7871
rect 12716 7828 12768 7837
rect 4252 7760 4304 7812
rect 4712 7760 4764 7812
rect 2688 7692 2740 7744
rect 4436 7692 4488 7744
rect 4896 7692 4948 7744
rect 5908 7803 5960 7812
rect 5908 7769 5917 7803
rect 5917 7769 5951 7803
rect 5951 7769 5960 7803
rect 5908 7760 5960 7769
rect 6644 7760 6696 7812
rect 8300 7803 8352 7812
rect 8300 7769 8309 7803
rect 8309 7769 8343 7803
rect 8343 7769 8352 7803
rect 8300 7760 8352 7769
rect 8576 7760 8628 7812
rect 11060 7760 11112 7812
rect 7288 7692 7340 7744
rect 8116 7692 8168 7744
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 8484 7692 8536 7744
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 10508 7735 10560 7744
rect 10508 7701 10533 7735
rect 10533 7701 10560 7735
rect 10508 7692 10560 7701
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 4528 7488 4580 7540
rect 6644 7488 6696 7540
rect 4988 7352 5040 7404
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 5816 7420 5868 7472
rect 6276 7420 6328 7472
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 6552 7352 6604 7404
rect 7564 7352 7616 7404
rect 8944 7488 8996 7540
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 11152 7488 11204 7540
rect 8208 7420 8260 7472
rect 10508 7420 10560 7472
rect 11980 7420 12032 7472
rect 9680 7395 9732 7404
rect 9680 7361 9689 7395
rect 9689 7361 9723 7395
rect 9723 7361 9732 7395
rect 9680 7352 9732 7361
rect 11152 7352 11204 7404
rect 11244 7395 11296 7404
rect 11244 7361 11263 7395
rect 11263 7361 11296 7395
rect 11244 7352 11296 7361
rect 12072 7352 12124 7404
rect 5356 7327 5408 7336
rect 5356 7293 5365 7327
rect 5365 7293 5399 7327
rect 5399 7293 5408 7327
rect 5356 7284 5408 7293
rect 10324 7284 10376 7336
rect 12532 7327 12584 7336
rect 12532 7293 12541 7327
rect 12541 7293 12575 7327
rect 12575 7293 12584 7327
rect 12532 7284 12584 7293
rect 3884 7259 3936 7268
rect 3884 7225 3893 7259
rect 3893 7225 3927 7259
rect 3927 7225 3936 7259
rect 3884 7216 3936 7225
rect 9036 7216 9088 7268
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 4620 7148 4672 7200
rect 5356 7148 5408 7200
rect 11980 7148 12032 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 5356 6987 5408 6996
rect 5356 6953 5365 6987
rect 5365 6953 5399 6987
rect 5399 6953 5408 6987
rect 5356 6944 5408 6953
rect 5908 6944 5960 6996
rect 7288 6944 7340 6996
rect 8208 6944 8260 6996
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 9220 6944 9272 6996
rect 9404 6944 9456 6996
rect 10692 6944 10744 6996
rect 12532 6944 12584 6996
rect 2688 6808 2740 6860
rect 4988 6876 5040 6928
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 848 6740 900 6792
rect 1584 6740 1636 6792
rect 2596 6740 2648 6792
rect 3148 6740 3200 6792
rect 4712 6783 4764 6792
rect 4712 6749 4721 6783
rect 4721 6749 4755 6783
rect 4755 6749 4764 6783
rect 4712 6740 4764 6749
rect 5264 6740 5316 6792
rect 5816 6783 5868 6792
rect 5816 6749 5825 6783
rect 5825 6749 5859 6783
rect 5859 6749 5868 6783
rect 5816 6740 5868 6749
rect 6000 6783 6052 6792
rect 6000 6749 6009 6783
rect 6009 6749 6043 6783
rect 6043 6749 6052 6783
rect 6000 6740 6052 6749
rect 6184 6740 6236 6792
rect 6460 6783 6512 6792
rect 6460 6749 6469 6783
rect 6469 6749 6503 6783
rect 6503 6749 6512 6783
rect 6460 6740 6512 6749
rect 1492 6672 1544 6724
rect 4804 6672 4856 6724
rect 5724 6672 5776 6724
rect 8484 6715 8536 6724
rect 8484 6681 8511 6715
rect 8511 6681 8536 6715
rect 8484 6672 8536 6681
rect 8576 6672 8628 6724
rect 8760 6672 8812 6724
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 2872 6604 2924 6656
rect 4344 6647 4396 6656
rect 4344 6613 4353 6647
rect 4353 6613 4387 6647
rect 4387 6613 4396 6647
rect 4344 6604 4396 6613
rect 4988 6604 5040 6656
rect 7932 6604 7984 6656
rect 8852 6604 8904 6656
rect 12808 6672 12860 6724
rect 9404 6604 9456 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1492 6400 1544 6452
rect 2872 6332 2924 6384
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 2136 6239 2188 6248
rect 2136 6205 2145 6239
rect 2145 6205 2179 6239
rect 2179 6205 2188 6239
rect 2136 6196 2188 6205
rect 4712 6400 4764 6452
rect 6828 6400 6880 6452
rect 8760 6400 8812 6452
rect 8944 6400 8996 6452
rect 9588 6400 9640 6452
rect 10232 6400 10284 6452
rect 11152 6400 11204 6452
rect 4804 6332 4856 6384
rect 4344 6264 4396 6316
rect 4620 6264 4672 6316
rect 8116 6375 8168 6384
rect 8116 6341 8125 6375
rect 8125 6341 8159 6375
rect 8159 6341 8168 6375
rect 8116 6332 8168 6341
rect 8208 6332 8260 6384
rect 11244 6375 11296 6384
rect 11244 6341 11253 6375
rect 11253 6341 11287 6375
rect 11287 6341 11296 6375
rect 11244 6332 11296 6341
rect 12072 6375 12124 6384
rect 12072 6341 12081 6375
rect 12081 6341 12115 6375
rect 12115 6341 12124 6375
rect 12072 6332 12124 6341
rect 3976 6128 4028 6180
rect 5080 6196 5132 6248
rect 5448 6196 5500 6248
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6552 6307 6604 6316
rect 6552 6273 6565 6307
rect 6565 6273 6604 6307
rect 6552 6264 6604 6273
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 8300 6264 8352 6316
rect 8576 6264 8628 6316
rect 9680 6264 9732 6316
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 9496 6196 9548 6248
rect 12532 6264 12584 6316
rect 2872 6060 2924 6112
rect 5264 6060 5316 6112
rect 5356 6103 5408 6112
rect 5356 6069 5365 6103
rect 5365 6069 5399 6103
rect 5399 6069 5408 6103
rect 5356 6060 5408 6069
rect 5724 6060 5776 6112
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 7012 6060 7064 6112
rect 8944 6060 8996 6112
rect 10232 6103 10284 6112
rect 10232 6069 10241 6103
rect 10241 6069 10275 6103
rect 10275 6069 10284 6103
rect 10232 6060 10284 6069
rect 10876 6060 10928 6112
rect 11704 6060 11756 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2136 5856 2188 5908
rect 2504 5899 2556 5908
rect 2504 5865 2513 5899
rect 2513 5865 2547 5899
rect 2547 5865 2556 5899
rect 2504 5856 2556 5865
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 2872 5831 2924 5840
rect 2872 5797 2881 5831
rect 2881 5797 2915 5831
rect 2915 5797 2924 5831
rect 2872 5788 2924 5797
rect 4804 5788 4856 5840
rect 2780 5652 2832 5704
rect 4712 5695 4764 5704
rect 4712 5661 4721 5695
rect 4721 5661 4755 5695
rect 4755 5661 4764 5695
rect 4712 5652 4764 5661
rect 6460 5856 6512 5908
rect 6552 5899 6604 5908
rect 6552 5865 6561 5899
rect 6561 5865 6595 5899
rect 6595 5865 6604 5899
rect 6552 5856 6604 5865
rect 7196 5856 7248 5908
rect 8852 5856 8904 5908
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 8944 5856 8996 5865
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 11520 5856 11572 5908
rect 11704 5856 11756 5908
rect 5172 5788 5224 5840
rect 2688 5584 2740 5636
rect 2596 5516 2648 5568
rect 4160 5627 4212 5636
rect 4160 5593 4169 5627
rect 4169 5593 4203 5627
rect 4203 5593 4212 5627
rect 4160 5584 4212 5593
rect 5172 5695 5224 5704
rect 5172 5661 5182 5695
rect 5182 5661 5216 5695
rect 5216 5661 5224 5695
rect 5448 5788 5500 5840
rect 6092 5788 6144 5840
rect 7012 5831 7064 5840
rect 7012 5797 7021 5831
rect 7021 5797 7055 5831
rect 7055 5797 7064 5831
rect 7012 5788 7064 5797
rect 8484 5788 8536 5840
rect 9312 5788 9364 5840
rect 9588 5788 9640 5840
rect 10232 5788 10284 5840
rect 5172 5652 5224 5661
rect 6460 5720 6512 5772
rect 6000 5695 6052 5704
rect 6000 5661 6009 5695
rect 6009 5661 6043 5695
rect 6043 5661 6052 5695
rect 6000 5652 6052 5661
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6552 5652 6604 5704
rect 6644 5695 6696 5704
rect 6644 5661 6653 5695
rect 6653 5661 6687 5695
rect 6687 5661 6696 5695
rect 6644 5652 6696 5661
rect 3332 5559 3384 5568
rect 3332 5525 3341 5559
rect 3341 5525 3375 5559
rect 3375 5525 3384 5559
rect 3332 5516 3384 5525
rect 3700 5516 3752 5568
rect 4344 5516 4396 5568
rect 4804 5516 4856 5568
rect 5540 5516 5592 5568
rect 5632 5516 5684 5568
rect 6368 5516 6420 5568
rect 7196 5652 7248 5704
rect 8392 5652 8444 5704
rect 8484 5695 8536 5704
rect 8484 5661 8493 5695
rect 8493 5661 8527 5695
rect 8527 5661 8536 5695
rect 8484 5652 8536 5661
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 9220 5652 9272 5704
rect 11244 5720 11296 5772
rect 9496 5652 9548 5704
rect 8116 5584 8168 5636
rect 8668 5584 8720 5636
rect 10048 5584 10100 5636
rect 8484 5559 8536 5568
rect 8484 5525 8493 5559
rect 8493 5525 8527 5559
rect 8527 5525 8536 5559
rect 8484 5516 8536 5525
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 9404 5516 9456 5568
rect 10784 5584 10836 5636
rect 11060 5584 11112 5636
rect 12808 5584 12860 5636
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 3792 5244 3844 5296
rect 4620 5312 4672 5364
rect 4712 5312 4764 5364
rect 4896 5312 4948 5364
rect 5356 5312 5408 5364
rect 6552 5312 6604 5364
rect 7196 5312 7248 5364
rect 11520 5355 11572 5364
rect 11520 5321 11529 5355
rect 11529 5321 11563 5355
rect 11563 5321 11572 5355
rect 11520 5312 11572 5321
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 5632 5244 5684 5296
rect 8668 5287 8720 5296
rect 8668 5253 8677 5287
rect 8677 5253 8711 5287
rect 8711 5253 8720 5287
rect 8668 5244 8720 5253
rect 9496 5287 9548 5296
rect 9496 5253 9505 5287
rect 9505 5253 9539 5287
rect 9539 5253 9548 5287
rect 9496 5244 9548 5253
rect 11336 5244 11388 5296
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 5264 5083 5316 5092
rect 5264 5049 5273 5083
rect 5273 5049 5307 5083
rect 5307 5049 5316 5083
rect 5264 5040 5316 5049
rect 9312 5219 9364 5228
rect 9312 5185 9321 5219
rect 9321 5185 9355 5219
rect 9355 5185 9364 5219
rect 9312 5176 9364 5185
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 10968 5176 11020 5228
rect 10232 5108 10284 5160
rect 11152 5108 11204 5160
rect 11980 5219 12032 5228
rect 11980 5185 11989 5219
rect 11989 5185 12023 5219
rect 12023 5185 12032 5219
rect 11980 5176 12032 5185
rect 12624 5176 12676 5228
rect 4068 4972 4120 5024
rect 4712 4972 4764 5024
rect 5172 5015 5224 5024
rect 5172 4981 5196 5015
rect 5196 4981 5224 5015
rect 5172 4972 5224 4981
rect 5632 5015 5684 5024
rect 5632 4981 5641 5015
rect 5641 4981 5675 5015
rect 5675 4981 5684 5015
rect 5632 4972 5684 4981
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 6828 4972 6880 5024
rect 8484 4972 8536 5024
rect 9680 4972 9732 5024
rect 12348 5015 12400 5024
rect 12348 4981 12357 5015
rect 12357 4981 12391 5015
rect 12391 4981 12400 5015
rect 12348 4972 12400 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2136 4768 2188 4820
rect 3332 4768 3384 4820
rect 3792 4768 3844 4820
rect 5356 4768 5408 4820
rect 6644 4768 6696 4820
rect 10048 4768 10100 4820
rect 3700 4700 3752 4752
rect 6460 4700 6512 4752
rect 10968 4768 11020 4820
rect 4712 4632 4764 4684
rect 3148 4564 3200 4616
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 7840 4632 7892 4684
rect 9680 4675 9732 4684
rect 9680 4641 9689 4675
rect 9689 4641 9723 4675
rect 9723 4641 9732 4675
rect 9680 4632 9732 4641
rect 2412 4496 2464 4548
rect 4068 4496 4120 4548
rect 6000 4496 6052 4548
rect 6184 4539 6236 4548
rect 6184 4505 6193 4539
rect 6193 4505 6227 4539
rect 6227 4505 6236 4539
rect 6184 4496 6236 4505
rect 7840 4539 7892 4548
rect 7840 4505 7849 4539
rect 7849 4505 7883 4539
rect 7883 4505 7892 4539
rect 7840 4496 7892 4505
rect 8024 4539 8076 4548
rect 8024 4505 8033 4539
rect 8033 4505 8067 4539
rect 8067 4505 8076 4539
rect 10784 4564 10836 4616
rect 11244 4564 11296 4616
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 12348 4607 12400 4616
rect 12348 4573 12349 4607
rect 12349 4573 12383 4607
rect 12383 4573 12400 4607
rect 12348 4564 12400 4573
rect 8024 4496 8076 4505
rect 9588 4496 9640 4548
rect 5264 4428 5316 4480
rect 6460 4428 6512 4480
rect 8116 4428 8168 4480
rect 8300 4471 8352 4480
rect 8300 4437 8309 4471
rect 8309 4437 8343 4471
rect 8343 4437 8352 4471
rect 8300 4428 8352 4437
rect 9312 4428 9364 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 3700 4224 3752 4276
rect 7840 4224 7892 4276
rect 7932 4224 7984 4276
rect 5724 4156 5776 4208
rect 9036 4224 9088 4276
rect 5632 4088 5684 4140
rect 5816 4088 5868 4140
rect 6184 4131 6236 4140
rect 6184 4097 6193 4131
rect 6193 4097 6227 4131
rect 6227 4097 6236 4131
rect 6184 4088 6236 4097
rect 6828 4088 6880 4140
rect 2780 4020 2832 4072
rect 4804 4020 4856 4072
rect 5356 4063 5408 4072
rect 5356 4029 5365 4063
rect 5365 4029 5399 4063
rect 5399 4029 5408 4063
rect 5356 4020 5408 4029
rect 8300 4020 8352 4072
rect 10232 4088 10284 4140
rect 9404 4020 9456 4072
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 12348 4088 12400 4140
rect 5908 3995 5960 4004
rect 5908 3961 5917 3995
rect 5917 3961 5951 3995
rect 5951 3961 5960 3995
rect 5908 3952 5960 3961
rect 8576 3952 8628 4004
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 7932 3927 7984 3936
rect 7932 3893 7941 3927
rect 7941 3893 7975 3927
rect 7975 3893 7984 3927
rect 7932 3884 7984 3893
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 4804 3680 4856 3732
rect 5356 3680 5408 3732
rect 6460 3723 6512 3732
rect 6460 3689 6469 3723
rect 6469 3689 6503 3723
rect 6503 3689 6512 3723
rect 6460 3680 6512 3689
rect 8760 3680 8812 3732
rect 8944 3680 8996 3732
rect 10232 3680 10284 3732
rect 12624 3680 12676 3732
rect 4620 3612 4672 3664
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 5908 3544 5960 3596
rect 6000 3587 6052 3596
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 6000 3544 6052 3553
rect 4804 3476 4856 3528
rect 5356 3519 5408 3528
rect 5356 3485 5365 3519
rect 5365 3485 5399 3519
rect 5399 3485 5408 3519
rect 5356 3476 5408 3485
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 8024 3544 8076 3596
rect 8944 3587 8996 3596
rect 8944 3553 8953 3587
rect 8953 3553 8987 3587
rect 8987 3553 8996 3587
rect 8944 3544 8996 3553
rect 9588 3544 9640 3596
rect 6184 3476 6236 3528
rect 6552 3519 6604 3528
rect 6552 3485 6561 3519
rect 6561 3485 6595 3519
rect 6595 3485 6604 3519
rect 6552 3476 6604 3485
rect 6644 3519 6696 3528
rect 6644 3485 6653 3519
rect 6653 3485 6687 3519
rect 6687 3485 6696 3519
rect 6644 3476 6696 3485
rect 6828 3519 6880 3528
rect 6828 3485 6837 3519
rect 6837 3485 6871 3519
rect 6871 3485 6880 3519
rect 6828 3476 6880 3485
rect 6920 3519 6972 3528
rect 6920 3485 6929 3519
rect 6929 3485 6963 3519
rect 6963 3485 6972 3519
rect 6920 3476 6972 3485
rect 7196 3476 7248 3528
rect 8300 3476 8352 3528
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 12992 3519 13044 3528
rect 12992 3485 13001 3519
rect 13001 3485 13035 3519
rect 13035 3485 13044 3519
rect 12992 3476 13044 3485
rect 5816 3340 5868 3392
rect 6644 3340 6696 3392
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 8576 3340 8628 3392
rect 10508 3408 10560 3460
rect 10232 3340 10284 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5356 3136 5408 3188
rect 8024 3136 8076 3188
rect 4620 3068 4672 3120
rect 6920 3068 6972 3120
rect 8576 3068 8628 3120
rect 9588 3068 9640 3120
rect 6000 3043 6052 3052
rect 6000 3009 6009 3043
rect 6009 3009 6043 3043
rect 6043 3009 6052 3043
rect 6000 3000 6052 3009
rect 6184 3043 6236 3052
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 6460 3000 6512 3052
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7564 3000 7616 3052
rect 7012 2932 7064 2984
rect 7932 2932 7984 2984
rect 6552 2907 6604 2916
rect 6552 2873 6561 2907
rect 6561 2873 6595 2907
rect 6595 2873 6604 2907
rect 6552 2864 6604 2873
rect 5816 2839 5868 2848
rect 5816 2805 5825 2839
rect 5825 2805 5859 2839
rect 5859 2805 5868 2839
rect 5816 2796 5868 2805
rect 7104 2796 7156 2848
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 5448 2592 5500 2644
rect 4804 2456 4856 2508
rect 7196 2592 7248 2644
rect 7472 2592 7524 2644
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 5816 2456 5868 2508
rect 8944 2456 8996 2508
rect 6736 2363 6788 2372
rect 6736 2329 6745 2363
rect 6745 2329 6779 2363
rect 6779 2329 6788 2363
rect 6736 2320 6788 2329
rect 7748 2320 7800 2372
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5170 15822 5226 16622
rect 5814 15822 5870 16622
rect 6458 15822 6514 16622
rect 7102 15822 7158 16622
rect 7746 15822 7802 16622
rect 8390 15822 8446 16622
rect 9034 15822 9090 16622
rect 9678 15822 9734 16622
rect 5184 14906 5212 15822
rect 5184 14878 5304 14906
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5276 13938 5304 14878
rect 5828 13938 5856 15822
rect 6472 13938 6500 15822
rect 7116 13938 7144 15822
rect 7760 13938 7788 15822
rect 8404 14006 8432 15822
rect 8392 14000 8444 14006
rect 8392 13942 8444 13948
rect 9048 13954 9076 15822
rect 9048 13938 9168 13954
rect 9692 13938 9720 15822
rect 5264 13932 5316 13938
rect 5264 13874 5316 13880
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7748 13932 7800 13938
rect 9048 13932 9180 13938
rect 9048 13926 9128 13932
rect 7748 13874 7800 13880
rect 9128 13874 9180 13880
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3608 13456 3660 13462
rect 3608 13398 3660 13404
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 3068 12442 3096 13194
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3056 12436 3108 12442
rect 3056 12378 3108 12384
rect 3528 12170 3556 12582
rect 3620 12442 3648 13398
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12850 3832 13126
rect 3792 12844 3844 12850
rect 3792 12786 3844 12792
rect 4172 12730 4200 13262
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12850 4292 13126
rect 4724 12850 4752 13738
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5816 13524 5868 13530
rect 5816 13466 5868 13472
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4712 12844 4764 12850
rect 4712 12786 4764 12792
rect 4528 12776 4580 12782
rect 4080 12702 4200 12730
rect 4342 12744 4398 12753
rect 4580 12724 4660 12730
rect 4528 12718 4660 12724
rect 4080 12442 4108 12702
rect 4540 12702 4660 12718
rect 4342 12679 4344 12688
rect 4396 12679 4398 12688
rect 4344 12650 4396 12656
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3608 12436 3660 12442
rect 3608 12378 3660 12384
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4526 12336 4582 12345
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 4344 12300 4396 12306
rect 4526 12271 4528 12280
rect 4344 12242 4396 12248
rect 4580 12271 4582 12280
rect 4528 12242 4580 12248
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3332 12096 3384 12102
rect 3332 12038 3384 12044
rect 3344 11694 3372 12038
rect 3528 11830 3556 12106
rect 3516 11824 3568 11830
rect 3516 11766 3568 11772
rect 3804 11762 3832 12242
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4172 11762 4200 12106
rect 4264 11898 4292 12174
rect 4356 11898 4384 12242
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 4448 12102 4476 12174
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4160 11756 4212 11762
rect 4160 11698 4212 11704
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3516 11008 3568 11014
rect 3516 10950 3568 10956
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 1688 10062 1716 10542
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2792 10130 2820 10406
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1676 10056 1728 10062
rect 1676 9998 1728 10004
rect 1504 9654 1532 9998
rect 1688 9654 1716 9998
rect 2044 9988 2096 9994
rect 2044 9930 2096 9936
rect 2056 9722 2084 9930
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 2320 9648 2372 9654
rect 2320 9590 2372 9596
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1872 8022 1900 8366
rect 2240 8090 2268 8774
rect 2332 8634 2360 9590
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2516 9042 2544 9386
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2608 8974 2636 9454
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 1860 8016 1912 8022
rect 1860 7958 1912 7964
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1596 6798 1624 7822
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 1584 6792 1636 6798
rect 1584 6734 1636 6740
rect 860 6361 888 6734
rect 1492 6724 1544 6730
rect 1492 6666 1544 6672
rect 1504 6458 1532 6666
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 846 6352 902 6361
rect 1504 6322 1532 6394
rect 1596 6322 1624 6734
rect 1872 6322 1900 7958
rect 2332 6914 2360 8570
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2424 8090 2452 8502
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2608 7886 2636 8774
rect 2792 8022 2820 10066
rect 2964 9716 3016 9722
rect 3068 9704 3096 10066
rect 3252 9722 3280 10542
rect 3528 10266 3556 10950
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3016 9676 3096 9704
rect 3240 9716 3292 9722
rect 2964 9658 3016 9664
rect 3240 9658 3292 9664
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 9450 2912 9522
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 9042 2912 9386
rect 2976 9110 3004 9658
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3068 9382 3096 9522
rect 3344 9382 3372 9862
rect 3528 9518 3556 10202
rect 3804 10130 3832 11698
rect 4080 11642 4108 11698
rect 3988 11614 4108 11642
rect 3988 11082 4016 11614
rect 4172 11540 4200 11698
rect 4632 11558 4660 12702
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 11626 4752 12650
rect 4816 11762 4844 13330
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5000 12209 5028 12922
rect 5078 12880 5134 12889
rect 5276 12850 5304 13330
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5644 12850 5672 13262
rect 5724 13252 5776 13258
rect 5724 13194 5776 13200
rect 5078 12815 5080 12824
rect 5132 12815 5134 12824
rect 5264 12844 5316 12850
rect 5080 12786 5132 12792
rect 5264 12786 5316 12792
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5080 12640 5132 12646
rect 5078 12608 5080 12617
rect 5172 12640 5224 12646
rect 5132 12608 5134 12617
rect 5172 12582 5224 12588
rect 5630 12608 5686 12617
rect 5078 12543 5134 12552
rect 5078 12472 5134 12481
rect 5078 12407 5134 12416
rect 5184 12434 5212 12582
rect 5630 12543 5686 12552
rect 5092 12306 5120 12407
rect 5184 12406 5304 12434
rect 5080 12300 5132 12306
rect 5080 12242 5132 12248
rect 4986 12200 5042 12209
rect 4986 12135 5042 12144
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4896 11892 4948 11898
rect 5276 11880 5304 12406
rect 5538 12200 5594 12209
rect 5538 12135 5594 12144
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 4896 11834 4948 11840
rect 5092 11852 5304 11880
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4080 11512 4200 11540
rect 4620 11552 4672 11558
rect 4080 11354 4108 11512
rect 4620 11494 4672 11500
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4724 11354 4752 11562
rect 4908 11354 4936 11834
rect 4988 11824 5040 11830
rect 4988 11766 5040 11772
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4908 11200 4936 11290
rect 4632 11172 4936 11200
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3896 10266 3924 10678
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3884 10260 3936 10266
rect 4632 10248 4660 11172
rect 5000 11150 5028 11766
rect 5092 11762 5120 11852
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5092 11218 5120 11698
rect 5172 11620 5224 11626
rect 5172 11562 5224 11568
rect 5184 11286 5212 11562
rect 5172 11280 5224 11286
rect 5172 11222 5224 11228
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4988 11144 5040 11150
rect 4816 11104 4988 11132
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4724 10266 4752 11018
rect 3884 10202 3936 10208
rect 4540 10220 4660 10248
rect 4712 10260 4764 10266
rect 3792 10124 3844 10130
rect 3792 10066 3844 10072
rect 4068 10056 4120 10062
rect 4120 10016 4292 10044
rect 4068 9998 4120 10004
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4172 9654 4200 9862
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 3332 9376 3384 9382
rect 3332 9318 3384 9324
rect 2964 9104 3016 9110
rect 2964 9046 3016 9052
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 8634 3648 8910
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 2872 8560 2924 8566
rect 2872 8502 2924 8508
rect 2884 8090 2912 8502
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2780 8016 2832 8022
rect 2780 7958 2832 7964
rect 3160 7886 3188 8230
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2332 6886 2452 6914
rect 846 6287 902 6296
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1872 5234 1900 6258
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2148 5914 2176 6190
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2148 4826 2176 5102
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2424 4554 2452 6886
rect 2700 6866 2728 7686
rect 2778 6896 2834 6905
rect 2688 6860 2740 6866
rect 2778 6831 2834 6840
rect 2688 6802 2740 6808
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 5914 2544 6598
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2608 5574 2636 6734
rect 2700 5642 2728 6802
rect 2792 5710 2820 6831
rect 3160 6798 3188 7822
rect 3896 7274 3924 9522
rect 4080 9160 4108 9590
rect 4264 9586 4292 10016
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4540 9382 4568 10220
rect 4712 10202 4764 10208
rect 4816 10146 4844 11104
rect 4988 11086 5040 11092
rect 5276 11014 5304 11698
rect 5368 11558 5396 12038
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5552 11132 5580 12135
rect 5644 11762 5672 12543
rect 5736 11898 5764 13194
rect 5828 12889 5856 13466
rect 5920 13394 5948 13670
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5814 12880 5870 12889
rect 5814 12815 5870 12824
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5644 11218 5672 11494
rect 5632 11212 5684 11218
rect 5632 11154 5684 11160
rect 5368 11104 5580 11132
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10674 5304 10950
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 4632 10118 4844 10146
rect 4632 9994 4660 10118
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4632 9586 4660 9930
rect 4620 9580 4672 9586
rect 4724 9568 4752 9998
rect 4816 9722 4844 9998
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4804 9580 4856 9586
rect 4724 9540 4804 9568
rect 4620 9522 4672 9528
rect 4804 9522 4856 9528
rect 4528 9376 4580 9382
rect 4528 9318 4580 9324
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4080 9132 4292 9160
rect 4264 8634 4292 9132
rect 4632 8974 4660 9522
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4724 8974 4752 9318
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 3988 8022 4016 8366
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 4264 7206 4292 7754
rect 4436 7744 4488 7750
rect 4632 7698 4660 8366
rect 4724 7818 4752 8774
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4436 7686 4488 7692
rect 4448 7290 4476 7686
rect 4540 7670 4660 7698
rect 4540 7546 4568 7670
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4448 7262 4660 7290
rect 4632 7206 4660 7262
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4620 7200 4672 7206
rect 4816 7154 4844 9522
rect 5264 8900 5316 8906
rect 5264 8842 5316 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 7750 4936 8366
rect 5000 8090 5028 8570
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4620 7142 4672 7148
rect 4724 7126 4844 7154
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4724 6798 4752 7126
rect 5000 6934 5028 7346
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 4712 6792 4764 6798
rect 4712 6734 4764 6740
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2884 6390 2912 6598
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2884 5846 2912 6054
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2688 5636 2740 5642
rect 2688 5578 2740 5584
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2412 4548 2464 4554
rect 2412 4490 2464 4496
rect 2792 4078 2820 5646
rect 3160 4622 3188 6734
rect 4344 6656 4396 6662
rect 4344 6598 4396 6604
rect 4356 6322 4384 6598
rect 4724 6458 4752 6734
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4712 6452 4764 6458
rect 4712 6394 4764 6400
rect 4816 6390 4844 6666
rect 5000 6662 5028 6870
rect 5276 6798 5304 8842
rect 5368 8242 5396 11104
rect 5448 11008 5500 11014
rect 5448 10950 5500 10956
rect 5460 10062 5488 10950
rect 5736 10674 5764 11834
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5552 10062 5580 10610
rect 5736 10062 5764 10610
rect 5828 10606 5856 12815
rect 5920 12322 5948 13330
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6288 12442 6316 13126
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 5920 12306 6132 12322
rect 5908 12300 6132 12306
rect 5960 12294 6132 12300
rect 5908 12242 5960 12248
rect 6104 12186 6132 12294
rect 6104 12158 6316 12186
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5920 11830 5948 12038
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5920 10742 5948 10950
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5448 10056 5500 10062
rect 5448 9998 5500 10004
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5724 10056 5776 10062
rect 5724 9998 5776 10004
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5552 9586 5580 9862
rect 5920 9654 5948 9930
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 5448 9512 5500 9518
rect 5500 9460 5580 9466
rect 5448 9454 5580 9460
rect 5460 9438 5580 9454
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8430 5488 8910
rect 5552 8498 5580 9438
rect 6104 9178 6132 9522
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5448 8424 5500 8430
rect 5448 8366 5500 8372
rect 5552 8294 5580 8434
rect 5540 8288 5592 8294
rect 5368 8214 5488 8242
rect 5540 8230 5592 8236
rect 5460 8106 5488 8214
rect 5356 8084 5408 8090
rect 5460 8078 5580 8106
rect 5356 8026 5408 8032
rect 5368 7342 5396 8026
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 7002 5396 7142
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4804 6384 4856 6390
rect 4804 6326 4856 6332
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4620 6316 4672 6322
rect 4620 6258 4672 6264
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5914 4016 6122
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3700 5568 3752 5574
rect 3700 5510 3752 5516
rect 3344 4826 3372 5510
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3712 4758 3740 5510
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3804 4826 3832 5238
rect 3988 5216 4016 5850
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4068 5228 4120 5234
rect 3988 5188 4068 5216
rect 4068 5170 4120 5176
rect 4172 5114 4200 5578
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4356 5234 4384 5510
rect 4632 5370 4660 6258
rect 4816 5846 4844 6326
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 5448 6248 5500 6254
rect 5448 6190 5500 6196
rect 4804 5840 4856 5846
rect 4710 5808 4766 5817
rect 4804 5782 4856 5788
rect 4710 5743 4766 5752
rect 4724 5710 4752 5743
rect 4712 5704 4764 5710
rect 5092 5692 5120 6190
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5170 5944 5226 5953
rect 5170 5879 5226 5888
rect 5184 5846 5212 5879
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 5172 5704 5224 5710
rect 5092 5664 5172 5692
rect 4712 5646 4764 5652
rect 5172 5646 5224 5652
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4724 5114 4752 5306
rect 4080 5086 4200 5114
rect 4632 5086 4752 5114
rect 4080 5030 4108 5086
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3700 4752 3752 4758
rect 3700 4694 3752 4700
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3712 4282 3740 4694
rect 4080 4554 4108 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3670 4660 5086
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4690 4752 4966
rect 4712 4684 4764 4690
rect 4712 4626 4764 4632
rect 4816 4622 4844 5510
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4908 4622 4936 5306
rect 5276 5098 5304 6054
rect 5368 5370 5396 6054
rect 5460 5846 5488 6190
rect 5448 5840 5500 5846
rect 5448 5782 5500 5788
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5264 5092 5316 5098
rect 5264 5034 5316 5040
rect 5172 5024 5224 5030
rect 5172 4966 5224 4972
rect 5184 4690 5212 4966
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3738 4844 4014
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4632 3126 4660 3606
rect 5276 3602 5304 4422
rect 5368 4078 5396 4762
rect 5356 4072 5408 4078
rect 5356 4014 5408 4020
rect 5368 3738 5396 4014
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 5356 3528 5408 3534
rect 5356 3470 5408 3476
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4816 2514 4844 3470
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5368 3194 5396 3470
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5460 2650 5488 5782
rect 5552 5692 5580 8078
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 6905 5672 7346
rect 5630 6896 5686 6905
rect 5630 6831 5686 6840
rect 5828 6798 5856 7414
rect 5920 7002 5948 7754
rect 6012 7410 6040 8026
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6012 6798 6040 7346
rect 6196 6798 6224 11698
rect 6288 11082 6316 12158
rect 6380 11626 6408 12650
rect 6472 11694 6500 13398
rect 6656 13326 6684 13738
rect 6736 13728 6788 13734
rect 6736 13670 6788 13676
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 6748 13530 6776 13670
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6564 12889 6592 13262
rect 6550 12880 6606 12889
rect 6550 12815 6552 12824
rect 6604 12815 6606 12824
rect 6552 12786 6604 12792
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6564 10674 6592 12786
rect 6656 11762 6684 13262
rect 6748 12646 6776 13466
rect 7012 13388 7064 13394
rect 7012 13330 7064 13336
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6826 13016 6882 13025
rect 6932 12986 6960 13126
rect 6826 12951 6882 12960
rect 6920 12980 6972 12986
rect 6840 12782 6868 12951
rect 6920 12922 6972 12928
rect 7024 12850 7052 13330
rect 7208 13326 7236 13670
rect 8312 13530 8340 13806
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 7208 12986 7236 13262
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6736 12640 6788 12646
rect 6736 12582 6788 12588
rect 6840 12238 6868 12718
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12481 6960 12582
rect 6918 12472 6974 12481
rect 7024 12442 7052 12786
rect 7484 12782 7512 13126
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7472 12776 7524 12782
rect 7378 12744 7434 12753
rect 7472 12718 7524 12724
rect 7378 12679 7380 12688
rect 7432 12679 7434 12688
rect 7380 12650 7432 12656
rect 6918 12407 6974 12416
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7484 12238 7512 12718
rect 7668 12617 7696 12786
rect 7654 12608 7710 12617
rect 7654 12543 7710 12552
rect 7760 12345 7788 12786
rect 7746 12336 7802 12345
rect 7852 12306 7880 13126
rect 7746 12271 7802 12280
rect 7840 12300 7892 12306
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 6656 10266 6684 10406
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6656 10062 6684 10202
rect 6748 10062 6776 10406
rect 7300 10062 7328 10406
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7104 9988 7156 9994
rect 7104 9930 7156 9936
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9654 6960 9862
rect 7116 9722 7144 9930
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7288 9920 7340 9926
rect 7288 9862 7340 9868
rect 7208 9722 7236 9862
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7196 9716 7248 9722
rect 7196 9658 7248 9664
rect 6920 9648 6972 9654
rect 6458 9616 6514 9625
rect 6920 9590 6972 9596
rect 7300 9586 7328 9862
rect 7392 9586 7420 10542
rect 7484 9926 7512 10610
rect 7760 10062 7788 12271
rect 7840 12242 7892 12248
rect 8128 12238 8156 13194
rect 8220 13025 8248 13262
rect 8206 13016 8262 13025
rect 8206 12951 8262 12960
rect 9416 12850 9444 13806
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9508 13326 9536 13670
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12918 9536 13262
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12986 9720 13126
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9586 12880 9642 12889
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 9404 12844 9456 12850
rect 9784 12866 9812 13738
rect 9876 13462 9904 13738
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9642 12838 9812 12866
rect 9876 12850 9904 13398
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 9968 12986 9996 13330
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10060 12850 10088 13194
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 9586 12815 9642 12824
rect 9404 12786 9456 12792
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8312 12374 8340 12718
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8300 12368 8352 12374
rect 8300 12310 8352 12316
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 7944 11762 7972 12038
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 7944 11218 7972 11698
rect 8404 11694 8432 12650
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8496 11830 8524 12242
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8588 11694 8616 12174
rect 8864 11762 8892 12786
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9496 12640 9548 12646
rect 9496 12582 9548 12588
rect 9128 12368 9180 12374
rect 9128 12310 9180 12316
rect 9140 12238 9168 12310
rect 9232 12238 9260 12582
rect 9508 12238 9536 12582
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 9128 12096 9180 12102
rect 9128 12038 9180 12044
rect 9232 12050 9260 12174
rect 9496 12096 9548 12102
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8404 11150 8432 11630
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8036 10674 8064 10950
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8036 10130 8064 10610
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8128 10062 8156 10406
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7472 9920 7524 9926
rect 7472 9862 7524 9868
rect 6458 9551 6514 9560
rect 6828 9580 6880 9586
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6288 8974 6316 9318
rect 6276 8968 6328 8974
rect 6276 8910 6328 8916
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 6288 7478 6316 7890
rect 6276 7472 6328 7478
rect 6276 7414 6328 7420
rect 6472 6798 6500 9551
rect 6828 9522 6880 9528
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 6656 8974 6684 9454
rect 6840 9178 6868 9522
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6564 7410 6592 8502
rect 6644 7812 6696 7818
rect 6644 7754 6696 7760
rect 6656 7546 6684 7754
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 6460 6792 6512 6798
rect 6460 6734 6512 6740
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5736 6118 5764 6666
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 5736 5817 5764 6054
rect 6012 5953 6040 6054
rect 5998 5944 6054 5953
rect 5998 5879 6054 5888
rect 5722 5808 5778 5817
rect 5722 5743 5778 5752
rect 6012 5710 6040 5879
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 6104 5710 6132 5782
rect 6000 5704 6052 5710
rect 5552 5664 5764 5692
rect 5540 5568 5592 5574
rect 5632 5568 5684 5574
rect 5540 5510 5592 5516
rect 5630 5536 5632 5545
rect 5684 5536 5686 5545
rect 5552 5386 5580 5510
rect 5630 5471 5686 5480
rect 5552 5358 5672 5386
rect 5644 5302 5672 5358
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4146 5672 4966
rect 5736 4214 5764 5664
rect 6000 5646 6052 5652
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6380 5574 6408 6258
rect 6564 5914 6592 6258
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6472 5778 6500 5850
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6368 5568 6420 5574
rect 6368 5510 6420 5516
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4554 6040 4966
rect 6472 4758 6500 5714
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6564 5545 6592 5646
rect 6550 5536 6606 5545
rect 6550 5471 6606 5480
rect 6564 5370 6592 5471
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6656 4826 6684 5646
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6460 4752 6512 4758
rect 6460 4694 6512 4700
rect 6000 4548 6052 4554
rect 6000 4490 6052 4496
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 6196 4146 6224 4490
rect 6460 4480 6512 4486
rect 6460 4422 6512 4428
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 6184 4140 6236 4146
rect 6184 4082 6236 4088
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3534 5580 3878
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5828 3398 5856 4082
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5920 3602 5948 3946
rect 6472 3738 6500 4422
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6000 3596 6052 3602
rect 6000 3538 6052 3544
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5828 2854 5856 3334
rect 6012 3058 6040 3538
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6644 3528 6696 3534
rect 6644 3470 6696 3476
rect 6196 3058 6224 3470
rect 6000 3052 6052 3058
rect 6000 2994 6052 3000
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1306 5304 2382
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 5828 800 5856 2450
rect 6472 800 6500 2994
rect 6564 2922 6592 3470
rect 6656 3398 6684 3470
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6748 2378 6776 8774
rect 6840 6458 6868 9114
rect 7196 9104 7248 9110
rect 7196 9046 7248 9052
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6840 5030 6868 6258
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 7024 5846 7052 6054
rect 7208 5914 7236 9046
rect 7760 8090 7788 9998
rect 8404 9636 8432 11086
rect 8496 10742 8524 11494
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 8404 9608 8524 9636
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8404 9042 8432 9318
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 8496 7886 8524 9608
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8588 7818 8616 11630
rect 8944 11552 8996 11558
rect 8944 11494 8996 11500
rect 8956 10674 8984 11494
rect 9048 10674 9076 12038
rect 9140 11762 9168 12038
rect 9232 12022 9352 12050
rect 9496 12038 9548 12044
rect 9324 11762 9352 12022
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8760 10192 8812 10198
rect 8760 10134 8812 10140
rect 8772 9450 8800 10134
rect 8864 9722 8892 10542
rect 8956 10062 8984 10610
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 9048 9994 9076 10610
rect 9036 9988 9088 9994
rect 9036 9930 9088 9936
rect 8852 9716 8904 9722
rect 8852 9658 8904 9664
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8576 7812 8628 7818
rect 8576 7754 8628 7760
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 7300 7002 7328 7686
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 5370 7236 5646
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6840 3534 6868 4082
rect 7208 3534 7236 5306
rect 6828 3528 6880 3534
rect 6828 3470 6880 3476
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 6932 3126 6960 3470
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7024 2990 7052 3334
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 7116 800 7144 2790
rect 7208 2650 7236 3470
rect 7576 3058 7604 7346
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7852 4554 7880 4626
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7852 4282 7880 4490
rect 7944 4282 7972 6598
rect 8128 6390 8156 7686
rect 8220 7478 8248 7686
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8312 7002 8340 7754
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8220 6390 8248 6938
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8208 6384 8260 6390
rect 8208 6326 8260 6332
rect 8128 5642 8156 6326
rect 8312 6322 8340 6938
rect 8496 6730 8524 7686
rect 8588 6730 8616 7754
rect 8956 7546 8984 7822
rect 9140 7732 9168 11698
rect 9508 11694 9536 12038
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9508 11150 9536 11630
rect 9692 11150 9720 11698
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9232 9994 9260 10678
rect 9508 10674 9536 10950
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9324 9586 9352 10610
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 9580 9364 9586
rect 9312 9522 9364 9528
rect 9220 9444 9272 9450
rect 9220 9386 9272 9392
rect 9232 8974 9260 9386
rect 9416 9178 9444 10542
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10198 9628 10406
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9692 10062 9720 10610
rect 9784 10062 9812 12838
rect 9864 12844 9916 12850
rect 9864 12786 9916 12792
rect 10048 12844 10100 12850
rect 10048 12786 10100 12792
rect 9876 12238 9904 12786
rect 9968 12294 10180 12322
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9968 12170 9996 12294
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 12164 10008 12170
rect 9956 12106 10008 12112
rect 10060 12102 10088 12174
rect 10152 12170 10180 12294
rect 10428 12238 10456 13126
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10612 12238 10640 12582
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 10888 11694 10916 12174
rect 11072 11762 11100 12174
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11150 10916 11630
rect 11072 11354 11100 11698
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11256 11218 11284 12786
rect 11334 12608 11390 12617
rect 11334 12543 11390 12552
rect 11348 12442 11376 12543
rect 11336 12436 11388 12442
rect 11336 12378 11388 12384
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11808 11898 11836 12174
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10606 10364 10950
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9692 9722 9720 9998
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9772 9376 9824 9382
rect 9876 9364 9904 10406
rect 10244 9654 10272 10474
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 9824 9336 9904 9364
rect 9772 9318 9824 9324
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9876 8974 9904 9336
rect 9220 8968 9272 8974
rect 9220 8910 9272 8916
rect 9864 8968 9916 8974
rect 9864 8910 9916 8916
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9220 7744 9272 7750
rect 9140 7704 9220 7732
rect 9220 7686 9272 7692
rect 8944 7540 8996 7546
rect 8944 7482 8996 7488
rect 8956 6866 8984 7482
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8484 6724 8536 6730
rect 8404 6684 8484 6712
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8404 5710 8432 6684
rect 8484 6666 8536 6672
rect 8576 6724 8628 6730
rect 8576 6666 8628 6672
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8588 6610 8616 6666
rect 8496 6582 8616 6610
rect 8496 5846 8524 6582
rect 8772 6458 8800 6666
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8496 5710 8524 5782
rect 8588 5710 8616 6258
rect 8864 5914 8892 6598
rect 8956 6458 8984 6802
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8944 6112 8996 6118
rect 8944 6054 8996 6060
rect 8956 5914 8984 6054
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8496 5030 8524 5510
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8024 4548 8076 4554
rect 8024 4490 8076 4496
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7932 4276 7984 4282
rect 7932 4218 7984 4224
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7484 2650 7512 2994
rect 7944 2990 7972 3878
rect 8036 3602 8064 4490
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8128 3942 8156 4422
rect 8312 4078 8340 4422
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 8036 3194 8064 3538
rect 8312 3534 8340 4014
rect 8588 4010 8616 5646
rect 8668 5636 8720 5642
rect 8668 5578 8720 5584
rect 8680 5302 8708 5578
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 9048 4282 9076 7210
rect 9232 7002 9260 7686
rect 9416 7546 9444 7890
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9232 5710 9260 6938
rect 9416 6662 9444 6938
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9324 5574 9352 5782
rect 9508 5710 9536 6190
rect 9600 5846 9628 6394
rect 9692 6322 9720 7346
rect 10244 6458 10272 9590
rect 10336 9450 10364 10542
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10704 10062 10732 10406
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10612 9654 10640 9998
rect 10600 9648 10652 9654
rect 10600 9590 10652 9596
rect 10704 9586 10732 9998
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10324 9444 10376 9450
rect 10324 9386 10376 9392
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10336 7342 10364 8434
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9588 5840 9640 5846
rect 9588 5782 9640 5788
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9324 5234 9352 5510
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4486 9352 5170
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9036 4276 9088 4282
rect 9036 4218 9088 4224
rect 9416 4078 9444 5510
rect 9508 5302 9536 5646
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9600 5234 9628 5782
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4554 9628 5170
rect 9680 5024 9732 5030
rect 9680 4966 9732 4972
rect 9692 4690 9720 4966
rect 9968 4808 9996 5850
rect 10244 5846 10272 6054
rect 10232 5840 10284 5846
rect 10232 5782 10284 5788
rect 10428 5658 10456 8026
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10520 7478 10548 7686
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10704 7002 10732 7686
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10888 6322 10916 11086
rect 11256 10742 11284 11154
rect 11900 10810 11928 11698
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11992 10742 12020 10950
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11980 10736 12032 10742
rect 11980 10678 12032 10684
rect 12084 10198 12112 11698
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 10968 10056 11020 10062
rect 10968 9998 11020 10004
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 12164 10056 12216 10062
rect 12268 10044 12296 11494
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10606 12480 11018
rect 12544 10674 12572 11766
rect 12636 10742 12664 11834
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12728 11218 12756 11494
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12728 10674 12756 11154
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12820 10985 12848 11086
rect 12806 10976 12862 10985
rect 12806 10911 12862 10920
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12452 10266 12480 10542
rect 12532 10532 12584 10538
rect 12532 10474 12584 10480
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12348 10056 12400 10062
rect 12268 10016 12348 10044
rect 12164 9998 12216 10004
rect 12348 9998 12400 10004
rect 10980 9382 11008 9998
rect 11256 9586 11284 9998
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 10980 9178 11008 9318
rect 10968 9172 11020 9178
rect 10968 9114 11020 9120
rect 10980 8430 11008 9114
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 11072 7954 11100 8366
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11072 7546 11100 7754
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11164 7410 11192 7482
rect 11256 7410 11284 9522
rect 11992 8974 12020 9930
rect 12084 9722 12112 9930
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 9330 12112 9454
rect 12176 9450 12204 9998
rect 12452 9874 12480 10202
rect 12544 10130 12572 10474
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12532 10124 12584 10130
rect 12532 10066 12584 10072
rect 12360 9846 12480 9874
rect 12360 9568 12388 9846
rect 12544 9722 12572 10066
rect 12636 10062 12664 10406
rect 12728 10266 12756 10610
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12440 9586 12492 9592
rect 12360 9540 12440 9568
rect 12164 9444 12216 9450
rect 12164 9386 12216 9392
rect 12360 9330 12388 9540
rect 12440 9528 12492 9534
rect 12636 9518 12664 9998
rect 12820 9704 12848 10610
rect 12912 10305 12940 11086
rect 12898 10296 12954 10305
rect 12898 10231 12954 10240
rect 12728 9676 12848 9704
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12084 9302 12388 9330
rect 12636 9178 12664 9454
rect 12728 9382 12756 9676
rect 12990 9616 13046 9625
rect 12808 9580 12860 9586
rect 12990 9551 13046 9560
rect 12808 9522 12860 9528
rect 12820 9450 12848 9522
rect 12808 9444 12860 9450
rect 12808 9386 12860 9392
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12820 9178 12848 9386
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 13004 8974 13032 9551
rect 11980 8968 12032 8974
rect 12716 8968 12768 8974
rect 11980 8910 12032 8916
rect 12714 8936 12716 8945
rect 12992 8968 13044 8974
rect 12768 8936 12770 8945
rect 11992 8072 12020 8910
rect 12992 8910 13044 8916
rect 12714 8871 12770 8880
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12072 8084 12124 8090
rect 11992 8044 12072 8072
rect 11992 7478 12020 8044
rect 12072 8026 12124 8032
rect 11980 7472 12032 7478
rect 11980 7414 12032 7420
rect 11152 7404 11204 7410
rect 11152 7346 11204 7352
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 12072 7404 12124 7410
rect 12072 7346 12124 7352
rect 11164 6712 11192 7346
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11164 6684 11284 6712
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10888 6118 10916 6258
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10060 5642 10456 5658
rect 10048 5636 10456 5642
rect 10100 5630 10456 5636
rect 10048 5578 10100 5584
rect 10428 5574 10456 5630
rect 10784 5636 10836 5642
rect 11060 5636 11112 5642
rect 10836 5596 11060 5624
rect 10784 5578 10836 5584
rect 11060 5578 11112 5584
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10244 5166 10272 5510
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10980 4826 11008 5170
rect 11164 5166 11192 6394
rect 11256 6390 11284 6684
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11256 5896 11284 6326
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11716 5914 11744 6054
rect 11520 5908 11572 5914
rect 11256 5868 11376 5896
rect 11244 5772 11296 5778
rect 11244 5714 11296 5720
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 10048 4820 10100 4826
rect 9968 4780 10048 4808
rect 10048 4762 10100 4768
rect 10968 4820 11020 4826
rect 10968 4762 11020 4768
rect 9680 4684 9732 4690
rect 9680 4626 9732 4632
rect 11256 4622 11284 5714
rect 11348 5302 11376 5868
rect 11520 5850 11572 5856
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11532 5370 11560 5850
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11716 4622 11744 5850
rect 11992 5234 12020 7142
rect 12084 6390 12112 7346
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12544 7002 12572 7278
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 12544 6322 12572 6938
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12636 5234 12664 8434
rect 12728 7886 12756 8434
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12820 6730 12848 8298
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12820 5370 12848 5578
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 11980 5228 12032 5234
rect 11980 5170 12032 5176
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4622 12388 4966
rect 10784 4616 10836 4622
rect 10784 4558 10836 4564
rect 11244 4616 11296 4622
rect 11244 4558 11296 4564
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 12348 4616 12400 4622
rect 12348 4558 12400 4564
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 8576 4004 8628 4010
rect 8576 3946 8628 3952
rect 8588 3534 8616 3946
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8772 3738 8800 3878
rect 8956 3738 8984 3878
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9600 3602 9628 4490
rect 10796 4146 10824 4558
rect 12360 4146 12388 4558
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 10244 3738 10272 4082
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8588 3126 8616 3334
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7760 2378 7788 2790
rect 8956 2514 8984 3538
rect 9600 3126 9628 3538
rect 10244 3398 10272 3674
rect 10520 3466 10548 3878
rect 12636 3738 12664 5170
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12992 3528 13044 3534
rect 12990 3496 12992 3505
rect 13044 3496 13046 3505
rect 10508 3460 10560 3466
rect 12990 3431 13046 3440
rect 10508 3402 10560 3408
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
<< via2 >>
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4342 12708 4398 12744
rect 4342 12688 4344 12708
rect 4344 12688 4396 12708
rect 4396 12688 4398 12708
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4526 12300 4582 12336
rect 4526 12280 4528 12300
rect 4528 12280 4580 12300
rect 4580 12280 4582 12300
rect 846 6296 902 6352
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 5078 12844 5134 12880
rect 5078 12824 5080 12844
rect 5080 12824 5132 12844
rect 5132 12824 5134 12844
rect 5078 12588 5080 12608
rect 5080 12588 5132 12608
rect 5132 12588 5134 12608
rect 5078 12552 5134 12588
rect 5078 12416 5134 12472
rect 5630 12552 5686 12608
rect 4986 12144 5042 12200
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 5538 12144 5594 12200
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 2778 6840 2834 6896
rect 5814 12824 5870 12880
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4710 5752 4766 5808
rect 5170 5888 5226 5944
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 5630 6840 5686 6896
rect 6550 12844 6606 12880
rect 6550 12824 6552 12844
rect 6552 12824 6604 12844
rect 6604 12824 6606 12844
rect 6826 12960 6882 13016
rect 6918 12416 6974 12472
rect 7378 12708 7434 12744
rect 7378 12688 7380 12708
rect 7380 12688 7432 12708
rect 7432 12688 7434 12708
rect 7654 12552 7710 12608
rect 7746 12280 7802 12336
rect 6458 9560 6514 9616
rect 8206 12960 8262 13016
rect 9586 12824 9642 12880
rect 5998 5888 6054 5944
rect 5722 5752 5778 5808
rect 5630 5516 5632 5536
rect 5632 5516 5684 5536
rect 5684 5516 5686 5536
rect 5630 5480 5686 5516
rect 6550 5480 6606 5536
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 11334 12552 11390 12608
rect 12806 10920 12862 10976
rect 12898 10240 12954 10296
rect 12990 9560 13046 9616
rect 12714 8916 12716 8936
rect 12716 8916 12768 8936
rect 12768 8916 12770 8936
rect 12714 8880 12770 8916
rect 12990 3476 12992 3496
rect 12992 3476 13044 3496
rect 13044 3476 13046 3496
rect 12990 3440 13046 3476
<< metal3 >>
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 6821 13018 6887 13021
rect 8201 13018 8267 13021
rect 6821 13016 8267 13018
rect 6821 12960 6826 13016
rect 6882 12960 8206 13016
rect 8262 12960 8267 13016
rect 6821 12958 8267 12960
rect 6821 12955 6887 12958
rect 8201 12955 8267 12958
rect 5073 12882 5139 12885
rect 5809 12882 5875 12885
rect 5073 12880 5875 12882
rect 5073 12824 5078 12880
rect 5134 12824 5814 12880
rect 5870 12824 5875 12880
rect 5073 12822 5875 12824
rect 5073 12819 5139 12822
rect 5809 12819 5875 12822
rect 6545 12882 6611 12885
rect 9581 12882 9647 12885
rect 6545 12880 9647 12882
rect 6545 12824 6550 12880
rect 6606 12824 9586 12880
rect 9642 12824 9647 12880
rect 6545 12822 9647 12824
rect 6545 12819 6611 12822
rect 9581 12819 9647 12822
rect 4337 12746 4403 12749
rect 7373 12746 7439 12749
rect 4337 12744 7439 12746
rect 4337 12688 4342 12744
rect 4398 12688 7378 12744
rect 7434 12688 7439 12744
rect 4337 12686 7439 12688
rect 4337 12683 4403 12686
rect 7373 12683 7439 12686
rect 5073 12610 5139 12613
rect 5625 12610 5691 12613
rect 5073 12608 5691 12610
rect 5073 12552 5078 12608
rect 5134 12552 5630 12608
rect 5686 12552 5691 12608
rect 5073 12550 5691 12552
rect 5073 12547 5139 12550
rect 5625 12547 5691 12550
rect 7649 12610 7715 12613
rect 11329 12610 11395 12613
rect 7649 12608 11395 12610
rect 7649 12552 7654 12608
rect 7710 12552 11334 12608
rect 11390 12552 11395 12608
rect 7649 12550 11395 12552
rect 7649 12547 7715 12550
rect 11329 12547 11395 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 5073 12474 5139 12477
rect 6913 12474 6979 12477
rect 5073 12472 6979 12474
rect 5073 12416 5078 12472
rect 5134 12416 6918 12472
rect 6974 12416 6979 12472
rect 5073 12414 6979 12416
rect 5073 12411 5139 12414
rect 6913 12411 6979 12414
rect 4521 12338 4587 12341
rect 7741 12338 7807 12341
rect 4521 12336 7807 12338
rect 4521 12280 4526 12336
rect 4582 12280 7746 12336
rect 7802 12280 7807 12336
rect 4521 12278 7807 12280
rect 4521 12275 4587 12278
rect 7741 12275 7807 12278
rect 4981 12202 5047 12205
rect 5533 12202 5599 12205
rect 4981 12200 5599 12202
rect 4981 12144 4986 12200
rect 5042 12144 5538 12200
rect 5594 12144 5599 12200
rect 4981 12142 5599 12144
rect 4981 12139 5047 12142
rect 5533 12139 5599 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12801 10978 12867 10981
rect 13678 10978 14478 11008
rect 12801 10976 14478 10978
rect 12801 10920 12806 10976
rect 12862 10920 14478 10976
rect 12801 10918 14478 10920
rect 12801 10915 12867 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 13678 10888 14478 10918
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12893 10298 12959 10301
rect 13678 10298 14478 10328
rect 12893 10296 14478 10298
rect 12893 10240 12898 10296
rect 12954 10240 14478 10296
rect 12893 10238 14478 10240
rect 12893 10235 12959 10238
rect 13678 10208 14478 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 6453 9618 6519 9621
rect 0 9616 6519 9618
rect 0 9560 6458 9616
rect 6514 9560 6519 9616
rect 0 9558 6519 9560
rect 0 9528 800 9558
rect 6453 9555 6519 9558
rect 12985 9618 13051 9621
rect 13678 9618 14478 9648
rect 12985 9616 14478 9618
rect 12985 9560 12990 9616
rect 13046 9560 14478 9616
rect 12985 9558 14478 9560
rect 12985 9555 13051 9558
rect 13678 9528 14478 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12709 8938 12775 8941
rect 13678 8938 14478 8968
rect 12709 8936 14478 8938
rect 12709 8880 12714 8936
rect 12770 8880 14478 8936
rect 12709 8878 14478 8880
rect 12709 8875 12775 8878
rect 13678 8848 14478 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 2773 6898 2839 6901
rect 5625 6898 5691 6901
rect 2773 6896 5691 6898
rect 2773 6840 2778 6896
rect 2834 6840 5630 6896
rect 5686 6840 5691 6896
rect 2773 6838 5691 6840
rect 2773 6835 2839 6838
rect 5625 6835 5691 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 0 6128 800 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 5165 5946 5231 5949
rect 5993 5946 6059 5949
rect 5165 5944 6059 5946
rect 5165 5888 5170 5944
rect 5226 5888 5998 5944
rect 6054 5888 6059 5944
rect 5165 5886 6059 5888
rect 5165 5883 5231 5886
rect 5993 5883 6059 5886
rect 4705 5810 4771 5813
rect 5717 5810 5783 5813
rect 4705 5808 5783 5810
rect 4705 5752 4710 5808
rect 4766 5752 5722 5808
rect 5778 5752 5783 5808
rect 4705 5750 5783 5752
rect 4705 5747 4771 5750
rect 5717 5747 5783 5750
rect 5625 5538 5691 5541
rect 6545 5538 6611 5541
rect 5625 5536 6611 5538
rect 5625 5480 5630 5536
rect 5686 5480 6550 5536
rect 6606 5480 6611 5536
rect 5625 5478 6611 5480
rect 5625 5475 5691 5478
rect 6545 5475 6611 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12985 3498 13051 3501
rect 13678 3498 14478 3528
rect 12985 3496 14478 3498
rect 12985 3440 12990 3496
rect 13046 3440 14478 3496
rect 12985 3438 14478 3440
rect 12985 3435 13051 3438
rect 13678 3408 14478 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 13632 4528 14192
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 14176 5188 14192
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _176_
timestamp -25199
transform 1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp -25199
transform 1 0 11040 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _178_
timestamp -25199
transform 1 0 7452 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179_
timestamp -25199
transform 1 0 9108 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _180_
timestamp -25199
transform -1 0 9844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp -25199
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _182_
timestamp -25199
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _183_
timestamp -25199
transform 1 0 5796 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _184_
timestamp -25199
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp -25199
transform -1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _186_
timestamp -25199
transform 1 0 5612 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp -25199
transform -1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _188_
timestamp -25199
transform 1 0 6808 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _189_
timestamp -25199
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _190_
timestamp -25199
transform -1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _191_
timestamp -25199
transform -1 0 12512 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _192_
timestamp -25199
transform -1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _193_
timestamp -25199
transform -1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _194_
timestamp -25199
transform -1 0 8188 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _195_
timestamp -25199
transform -1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _196_
timestamp -25199
transform -1 0 6256 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _197_
timestamp -25199
transform -1 0 6992 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_1  _198_
timestamp -25199
transform -1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _199_
timestamp -25199
transform 1 0 4876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _200_
timestamp -25199
transform -1 0 6716 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _201_
timestamp -25199
transform -1 0 4048 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _202_
timestamp -25199
transform 1 0 3864 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _203_
timestamp -25199
transform 1 0 3680 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _204_
timestamp -25199
transform -1 0 6256 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _205_
timestamp -25199
transform 1 0 4692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _206_
timestamp -25199
transform -1 0 6072 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _207_
timestamp -25199
transform -1 0 5060 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _208_
timestamp -25199
transform -1 0 8648 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _209_
timestamp -25199
transform -1 0 7360 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _210_
timestamp -25199
transform 1 0 7728 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _211_
timestamp -25199
transform 1 0 6992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _212_
timestamp -25199
transform 1 0 7728 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _213_
timestamp -25199
transform 1 0 9384 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _214_
timestamp -25199
transform 1 0 8464 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _215_
timestamp -25199
transform -1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _216_
timestamp -25199
transform 1 0 10120 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _217_
timestamp -25199
transform 1 0 10028 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _218_
timestamp -25199
transform 1 0 12420 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _219_
timestamp -25199
transform 1 0 11316 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _220_
timestamp -25199
transform -1 0 11316 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _221_
timestamp -25199
transform -1 0 12880 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _222_
timestamp -25199
transform 1 0 12328 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _223_
timestamp -25199
transform -1 0 11316 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _224_
timestamp -25199
transform -1 0 12052 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _225_
timestamp -25199
transform -1 0 12604 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _226_
timestamp -25199
transform -1 0 12420 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _227_
timestamp -25199
transform -1 0 12144 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _228_
timestamp -25199
transform 1 0 11316 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _229_
timestamp -25199
transform 1 0 7360 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _230_
timestamp -25199
transform -1 0 4968 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _231_
timestamp -25199
transform -1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _232_
timestamp -25199
transform 1 0 4784 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _233_
timestamp -25199
transform -1 0 5060 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _234_
timestamp -25199
transform -1 0 5612 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _235_
timestamp -25199
transform 1 0 4600 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _236_
timestamp -25199
transform -1 0 6256 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _237_
timestamp -25199
transform 1 0 6900 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _238_
timestamp -25199
transform 1 0 5336 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _239_
timestamp -25199
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _240_
timestamp -25199
transform 1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp -25199
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _242_
timestamp -25199
transform -1 0 6348 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _243_
timestamp -25199
transform 1 0 6624 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _244_
timestamp -25199
transform 1 0 4968 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_1  _245_
timestamp -25199
transform -1 0 3680 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _246_
timestamp -25199
transform -1 0 4876 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _247_
timestamp -25199
transform 1 0 3036 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _248_
timestamp -25199
transform 1 0 3864 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _249_
timestamp -25199
transform -1 0 4692 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _250_
timestamp -25199
transform -1 0 5980 0 -1 4352
box -38 -48 1050 592
use sky130_fd_sc_hd__a21oi_1  _251_
timestamp -25199
transform -1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _252_
timestamp -25199
transform 1 0 5060 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _253_
timestamp -25199
transform 1 0 5060 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _254_
timestamp -25199
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _255_
timestamp -25199
transform 1 0 10580 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _256_
timestamp -25199
transform -1 0 11960 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _257_
timestamp -25199
transform 1 0 10304 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _258_
timestamp -25199
transform -1 0 10672 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _259_
timestamp -25199
transform 1 0 11500 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _260_
timestamp -25199
transform -1 0 10856 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _261_
timestamp -25199
transform -1 0 11316 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp -25199
transform 1 0 11500 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _263_
timestamp -25199
transform 1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _264_
timestamp -25199
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _265_
timestamp -25199
transform -1 0 9568 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _266_
timestamp -25199
transform 1 0 8648 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _267_
timestamp -25199
transform -1 0 8740 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _268_
timestamp -25199
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _269_
timestamp -25199
transform 1 0 7728 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _270_
timestamp -25199
transform -1 0 9568 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _271_
timestamp -25199
transform 1 0 8280 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _272_
timestamp -25199
transform 1 0 7636 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _273_
timestamp -25199
transform -1 0 6072 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _274_
timestamp -25199
transform -1 0 6256 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _275_
timestamp -25199
transform 1 0 4968 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _276_
timestamp -25199
transform -1 0 4968 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _277_
timestamp -25199
transform -1 0 5060 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _278_
timestamp -25199
transform 1 0 3864 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _279_
timestamp -25199
transform -1 0 3588 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _280_
timestamp -25199
transform -1 0 3128 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _281_
timestamp -25199
transform -1 0 2668 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _282_
timestamp -25199
transform 1 0 1472 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _283_
timestamp -25199
transform 1 0 1564 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _284_
timestamp -25199
transform -1 0 4048 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _285_
timestamp -25199
transform -1 0 3588 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _286_
timestamp -25199
transform 1 0 2484 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _287_
timestamp -25199
transform 1 0 1840 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _288_
timestamp -25199
transform 1 0 1380 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _289_
timestamp -25199
transform 1 0 2116 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _290_
timestamp -25199
transform -1 0 2944 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _291_
timestamp -25199
transform -1 0 4232 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _292_
timestamp -25199
transform 1 0 2944 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _293_
timestamp -25199
transform -1 0 2668 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _294_
timestamp -25199
transform -1 0 8740 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _295_
timestamp -25199
transform 1 0 7820 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _296_
timestamp -25199
transform -1 0 8556 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _297_
timestamp -25199
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _298_
timestamp -25199
transform 1 0 9936 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _299_
timestamp -25199
transform 1 0 8556 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _300_
timestamp -25199
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _301_
timestamp -25199
transform 1 0 5060 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _302_
timestamp -25199
transform 1 0 6164 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _303_
timestamp -25199
transform 1 0 5796 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _304_
timestamp -25199
transform 1 0 6348 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _305_
timestamp -25199
transform -1 0 4784 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _306_
timestamp -25199
transform 1 0 4508 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_2  _307_
timestamp -25199
transform 1 0 4784 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_1  _308_
timestamp -25199
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o22ai_1  _309_
timestamp -25199
transform 1 0 6532 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _310_
timestamp -25199
transform -1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _311_
timestamp -25199
transform -1 0 8556 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _312_
timestamp -25199
transform -1 0 8556 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _313_
timestamp -25199
transform -1 0 9568 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _314_
timestamp -25199
transform 1 0 9016 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _315_
timestamp -25199
transform 1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _316_
timestamp -25199
transform -1 0 10304 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _317_
timestamp -25199
transform -1 0 10948 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _318_
timestamp -25199
transform 1 0 10396 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _319_
timestamp -25199
transform -1 0 10396 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _320_
timestamp -25199
transform -1 0 9568 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _321_
timestamp -25199
transform -1 0 9476 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _322_
timestamp -25199
transform -1 0 9752 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _323_
timestamp -25199
transform 1 0 8556 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _324_
timestamp -25199
transform 1 0 7820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _325_
timestamp -25199
transform 1 0 6992 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _326_
timestamp -25199
transform -1 0 6992 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _327_
timestamp -25199
transform 1 0 5336 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _328_
timestamp -25199
transform -1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _329_
timestamp -25199
transform -1 0 7360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _330_
timestamp -25199
transform 1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_1  _331_
timestamp -25199
transform -1 0 9660 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or4b_4  _332_
timestamp -25199
transform -1 0 9292 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__and4bb_1  _333_
timestamp -25199
transform -1 0 8832 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__nand4b_1  _334_
timestamp -25199
transform -1 0 6256 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _335_
timestamp -25199
transform -1 0 6900 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _336_
timestamp -25199
transform 1 0 12696 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _337_
timestamp -25199
transform 1 0 12696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _338_
timestamp -25199
transform -1 0 12420 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _339_
timestamp -25199
transform 1 0 12696 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp -25199
transform -1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _341_
timestamp -25199
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp -25199
transform -1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _343_
timestamp -25199
transform 1 0 6624 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _344_
timestamp -25199
transform -1 0 6072 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _345_
timestamp -25199
transform -1 0 4324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _346_
timestamp -25199
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp -25199
transform 1 0 2852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _348_
timestamp -25199
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp -25199
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _350_
timestamp -25199
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _351_
timestamp -25199
transform -1 0 10672 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _352_
timestamp -25199
transform 1 0 6440 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _353_
timestamp -25199
transform 1 0 10764 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _354_
timestamp -25199
transform 1 0 11040 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _355_
timestamp -25199
transform 1 0 9568 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _356_
timestamp -25199
transform 1 0 10856 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _357_
timestamp -25199
transform 1 0 9384 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _358_
timestamp -25199
transform 1 0 8924 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _359_
timestamp -25199
transform 1 0 7636 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _360_
timestamp -25199
transform 1 0 5612 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _361_
timestamp -25199
transform 1 0 3956 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _362_
timestamp -25199
transform 1 0 1748 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _363_
timestamp -25199
transform -1 0 3588 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _364_
timestamp -25199
transform 1 0 1840 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _365_
timestamp -25199
transform 1 0 1840 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _366_
timestamp -25199
transform 1 0 1840 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _367_
timestamp -25199
transform -1 0 9936 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _368_
timestamp -25199
transform 1 0 8924 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 6440 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -25199
transform -1 0 5612 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -25199
transform 1 0 8372 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_2  clkload0
timestamp -25199
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  clone4
timestamp -25199
transform -1 0 5796 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout19
timestamp -25199
transform -1 0 2300 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout20
timestamp -25199
transform 1 0 9108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout21
timestamp -25199
transform -1 0 12696 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp -25199
transform 1 0 12144 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41
timestamp -25199
transform 1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp -25199
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp -25199
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636943256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -25199
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636943256
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp -25199
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp -25199
transform 1 0 12972 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636943256
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636943256
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636943256
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_39
timestamp -25199
transform 1 0 4692 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_45
timestamp -25199
transform 1 0 5244 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp -25199
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp -25199
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_70
timestamp -25199
transform 1 0 7544 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_74
timestamp -25199
transform 1 0 7912 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_96
timestamp 1636943256
transform 1 0 9936 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp -25199
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636943256
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp -25199
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129
timestamp -25199
transform 1 0 12972 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636943256
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636943256
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp -25199
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp -25199
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_35
timestamp -25199
transform 1 0 4324 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_66
timestamp -25199
transform 1 0 7176 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_74
timestamp -25199
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_80
timestamp -25199
transform 1 0 8464 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_105
timestamp 1636943256
transform 1 0 10764 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_117
timestamp -25199
transform 1 0 11868 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp -25199
transform 1 0 12604 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636943256
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636943256
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_27
timestamp -25199
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636943256
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp -25199
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_73
timestamp -25199
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_86
timestamp -25199
transform 1 0 9016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp -25199
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp -25199
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636943256
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_125
timestamp -25199
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp -25199
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp -25199
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp -25199
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_17
timestamp -25199
transform 1 0 2668 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp -25199
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_32
timestamp -25199
transform 1 0 4048 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_42
timestamp -25199
transform 1 0 4968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_48
timestamp -25199
transform 1 0 5520 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_54
timestamp -25199
transform 1 0 6072 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_62
timestamp -25199
transform 1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_70
timestamp -25199
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp -25199
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp -25199
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_118
timestamp -25199
transform 1 0 11960 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_123
timestamp -25199
transform 1 0 12420 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_129
timestamp -25199
transform 1 0 12972 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp -25199
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp -25199
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636943256
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636943256
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_81
timestamp -25199
transform 1 0 8556 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_119
timestamp -25199
transform 1 0 12052 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_129
timestamp -25199
transform 1 0 12972 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp -25199
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp -25199
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_68
timestamp -25199
transform 1 0 7360 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp -25199
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp -25199
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp -25199
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_29
timestamp -25199
transform 1 0 3772 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_37
timestamp -25199
transform 1 0 4508 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -25199
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_65
timestamp -25199
transform 1 0 7084 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_71
timestamp -25199
transform 1 0 7636 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp -25199
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp -25199
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp -25199
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_127
timestamp -25199
transform 1 0 12788 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_6
timestamp -25199
transform 1 0 1656 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_10
timestamp -25199
transform 1 0 2024 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_16
timestamp -25199
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_8_22
timestamp -25199
transform 1 0 3128 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_29
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp -25199
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp -25199
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_106
timestamp -25199
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_129
timestamp -25199
transform 1 0 12972 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636943256
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636943256
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp -25199
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_63
timestamp -25199
transform 1 0 6900 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_94
timestamp 1636943256
transform 1 0 9752 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp -25199
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp -25199
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_125
timestamp -25199
transform 1 0 12604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_129
timestamp -25199
transform 1 0 12972 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp -25199
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_7
timestamp -25199
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_15
timestamp -25199
transform 1 0 2484 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_22
timestamp -25199
transform 1 0 3128 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_70
timestamp -25199
transform 1 0 7544 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp -25199
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_92
timestamp -25199
transform 1 0 9568 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_129
timestamp -25199
transform 1 0 12972 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp -25199
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_7
timestamp -25199
transform 1 0 1748 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp -25199
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp -25199
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1636943256
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1636943256
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1636943256
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_93
timestamp -25199
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp -25199
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp -25199
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_113
timestamp -25199
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_119
timestamp -25199
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_129
timestamp -25199
transform 1 0 12972 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636943256
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp -25199
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp -25199
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp -25199
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_43
timestamp 1636943256
transform 1 0 5060 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_55
timestamp -25199
transform 1 0 6164 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_63
timestamp 1636943256
transform 1 0 6900 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_75
timestamp -25199
transform 1 0 8004 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp -25199
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp -25199
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_91
timestamp 1636943256
transform 1 0 9476 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_103
timestamp -25199
transform 1 0 10580 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_109
timestamp -25199
transform 1 0 11132 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_113
timestamp -25199
transform 1 0 11500 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_121
timestamp -25199
transform 1 0 12236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp -25199
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_35
timestamp -25199
transform 1 0 4324 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp -25199
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp -25199
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_69
timestamp -25199
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_77
timestamp -25199
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp -25199
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_100
timestamp -25199
transform 1 0 10304 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_107
timestamp -25199
transform 1 0 10948 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -25199
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_128
timestamp -25199
transform 1 0 12880 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp -25199
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_32
timestamp -25199
transform 1 0 4048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_52
timestamp -25199
transform 1 0 5888 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_68
timestamp -25199
transform 1 0 7360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp -25199
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_128
timestamp -25199
transform 1 0 12880 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp -25199
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636943256
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_39
timestamp -25199
transform 1 0 4692 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp -25199
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp -25199
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp -25199
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_64
timestamp -25199
transform 1 0 6992 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_72
timestamp -25199
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_79
timestamp -25199
transform 1 0 8372 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_94
timestamp -25199
transform 1 0 9752 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp -25199
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp -25199
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_128
timestamp -25199
transform 1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636943256
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636943256
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp -25199
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp -25199
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_43
timestamp -25199
transform 1 0 5060 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_49
timestamp -25199
transform 1 0 5612 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_54
timestamp 1636943256
transform 1 0 6072 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_66
timestamp -25199
transform 1 0 7176 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_74
timestamp -25199
transform 1 0 7912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp -25199
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_85
timestamp -25199
transform 1 0 8924 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp -25199
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_93
timestamp 1636943256
transform 1 0 9660 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_105
timestamp -25199
transform 1 0 10764 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_117
timestamp -25199
transform 1 0 11868 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636943256
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_15
timestamp -25199
transform 1 0 2484 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_36
timestamp -25199
transform 1 0 4416 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_40
timestamp -25199
transform 1 0 4784 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp -25199
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_60
timestamp 1636943256
transform 1 0 6624 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_72
timestamp -25199
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp -25199
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_85
timestamp -25199
transform 1 0 8924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636943256
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp -25199
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp -25199
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_125
timestamp -25199
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_129
timestamp -25199
transform 1 0 12972 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636943256
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_15
timestamp -25199
transform 1 0 2484 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp -25199
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_41
timestamp -25199
transform 1 0 4876 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp -25199
transform 1 0 6256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_60
timestamp -25199
transform 1 0 6624 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_64
timestamp -25199
transform 1 0 6992 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp -25199
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_95
timestamp -25199
transform 1 0 9844 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_117
timestamp 1636943256
transform 1 0 11868 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_129
timestamp -25199
transform 1 0 12972 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636943256
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_15
timestamp -25199
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_23
timestamp -25199
transform 1 0 3220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_79
timestamp -25199
transform 1 0 8372 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp -25199
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp -25199
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp -25199
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636943256
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp -25199
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_129
timestamp -25199
transform 1 0 12972 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1636943256
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1636943256
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp -25199
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp -25199
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_36
timestamp 1636943256
transform 1 0 4416 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_48
timestamp -25199
transform 1 0 5520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp -25199
transform 1 0 6716 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp -25199
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_85
timestamp -25199
transform 1 0 8924 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp -25199
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1636943256
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1636943256
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_121
timestamp -25199
transform 1 0 12236 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_129
timestamp -25199
transform 1 0 12972 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636943256
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636943256
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_27
timestamp -25199
transform 1 0 3588 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_29
timestamp 1636943256
transform 1 0 3772 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp -25199
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_48
timestamp -25199
transform 1 0 5520 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp -25199
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp -25199
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp -25199
transform 1 0 6808 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_69
timestamp -25199
transform 1 0 7452 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_82
timestamp -25199
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp -25199
transform 1 0 9568 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp -25199
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp -25199
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636943256
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp -25199
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp -25199
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -25199
transform 1 0 12788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp -25199
transform 1 0 5244 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -25199
transform -1 0 6164 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp -25199
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -25199
transform -1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp -25199
transform -1 0 6256 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -25199
transform -1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input8
timestamp -25199
transform -1 0 13064 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp -25199
transform 1 0 12512 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -25199
transform -1 0 12236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input11
timestamp -25199
transform 1 0 9752 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input12
timestamp -25199
transform 1 0 9292 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input13
timestamp -25199
transform 1 0 7820 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input14
timestamp -25199
transform 1 0 7176 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp -25199
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp -25199
transform -1 0 6808 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp -25199
transform -1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -25199
transform -1 0 7544 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_22
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_23
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_24
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_25
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_26
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_27
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_28
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_29
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 13340 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_30
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_31
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_32
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 13340 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_33
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 13340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_34
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 13340 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_35
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_36
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_37
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 13340 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_38
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_39
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_40
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 13340 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_41
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 13340 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_42
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_43
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer1
timestamp -25199
transform -1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp -25199
transform -1 0 6256 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp -25199
transform 1 0 4324 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer5
timestamp -25199
transform -1 0 12604 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  rebuffer6
timestamp -25199
transform -1 0 12788 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp -25199
transform 1 0 11040 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_44
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_45
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_48
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_49
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_50
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_51
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_52
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_53
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_54
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_55
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_56
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_57
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_58
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_59
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_60
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_61
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_62
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_63
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_64
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_65
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_66
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_67
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_68
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_69
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_70
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_71
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_72
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_73
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_74
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_75
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_76
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_77
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_78
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_79
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_80
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_81
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_82
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_83
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_84
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_85
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_86
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_87
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_88
timestamp -25199
transform 1 0 3680 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_89
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_90
timestamp -25199
transform 1 0 8832 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_91
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 14192 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 14192 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 out
port 3 nsew signal output
flabel metal3 s 13678 9528 14478 9648 0 FreeSans 480 0 0 0 psc[0]
port 4 nsew signal input
flabel metal2 s 5170 15822 5226 16622 0 FreeSans 224 90 0 0 psc[10]
port 5 nsew signal input
flabel metal2 s 5814 15822 5870 16622 0 FreeSans 224 90 0 0 psc[11]
port 6 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 psc[12]
port 7 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 psc[13]
port 8 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 psc[14]
port 9 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 psc[15]
port 10 nsew signal input
flabel metal3 s 13678 10208 14478 10328 0 FreeSans 480 0 0 0 psc[1]
port 11 nsew signal input
flabel metal3 s 13678 8848 14478 8968 0 FreeSans 480 0 0 0 psc[2]
port 12 nsew signal input
flabel metal3 s 13678 10888 14478 11008 0 FreeSans 480 0 0 0 psc[3]
port 13 nsew signal input
flabel metal2 s 9678 15822 9734 16622 0 FreeSans 224 90 0 0 psc[4]
port 14 nsew signal input
flabel metal2 s 9034 15822 9090 16622 0 FreeSans 224 90 0 0 psc[5]
port 15 nsew signal input
flabel metal2 s 7746 15822 7802 16622 0 FreeSans 224 90 0 0 psc[6]
port 16 nsew signal input
flabel metal2 s 7102 15822 7158 16622 0 FreeSans 224 90 0 0 psc[7]
port 17 nsew signal input
flabel metal2 s 8390 15822 8446 16622 0 FreeSans 224 90 0 0 psc[8]
port 18 nsew signal input
flabel metal2 s 6458 15822 6514 16622 0 FreeSans 224 90 0 0 psc[9]
port 19 nsew signal input
flabel metal3 s 13678 3408 14478 3528 0 FreeSans 480 0 0 0 rst
port 20 nsew signal input
rlabel metal1 7222 14144 7222 14144 0 VGND
rlabel metal1 7222 13600 7222 13600 0 VPWR
rlabel metal2 11086 8160 11086 8160 0 _000_
rlabel metal1 3450 9690 3450 9690 0 _001_
rlabel metal2 2438 8296 2438 8296 0 _002_
rlabel metal1 2254 5882 2254 5882 0 _003_
rlabel metal1 2116 4794 2116 4794 0 _004_
rlabel metal1 8786 2958 8786 2958 0 _005_
rlabel metal1 9098 3706 9098 3706 0 _006_
rlabel metal1 11030 6970 11030 6970 0 _007_
rlabel metal1 10074 5134 10074 5134 0 _008_
rlabel metal1 11132 5610 11132 5610 0 _009_
rlabel metal2 9706 4828 9706 4828 0 _010_
rlabel metal1 8556 6426 8556 6426 0 _011_
rlabel metal1 8096 7446 8096 7446 0 _012_
rlabel metal1 5750 6970 5750 6970 0 _013_
rlabel metal1 4508 7514 4508 7514 0 _014_
rlabel metal2 2070 9826 2070 9826 0 _015_
rlabel metal1 6808 8806 6808 8806 0 _016_
rlabel metal2 7774 2584 7774 2584 0 _017_
rlabel metal1 12565 7786 12565 7786 0 _018_
rlabel metal1 12703 6698 12703 6698 0 _019_
rlabel metal1 11638 4794 11638 4794 0 _020_
rlabel metal2 12834 5474 12834 5474 0 _021_
rlabel metal2 10810 4352 10810 4352 0 _022_
rlabel metal1 8786 5882 8786 5882 0 _023_
rlabel metal1 9391 7446 9391 7446 0 _024_
rlabel metal1 6716 7514 6716 7514 0 _025_
rlabel metal1 5711 8534 5711 8534 0 _026_
rlabel metal2 4186 9758 4186 9758 0 _027_
rlabel metal2 3910 10472 3910 10472 0 _028_
rlabel metal1 2944 8058 2944 8058 0 _029_
rlabel metal2 2898 6494 2898 6494 0 _030_
rlabel metal1 3864 4794 3864 4794 0 _031_
rlabel metal1 8648 3366 8648 3366 0 _032_
rlabel metal1 10495 3434 10495 3434 0 _033_
rlabel metal1 7544 13226 7544 13226 0 _034_
rlabel metal1 7314 12852 7314 12852 0 _035_
rlabel metal1 8142 12784 8142 12784 0 _036_
rlabel metal1 6992 12614 6992 12614 0 _037_
rlabel metal1 7406 12920 7406 12920 0 _038_
rlabel metal1 10212 13158 10212 13158 0 _039_
rlabel metal1 8050 12886 8050 12886 0 _040_
rlabel metal1 10672 12682 10672 12682 0 _041_
rlabel metal1 10534 12274 10534 12274 0 _042_
rlabel metal1 11408 12206 11408 12206 0 _043_
rlabel metal2 12742 10438 12742 10438 0 _044_
rlabel metal1 11408 11730 11408 11730 0 _045_
rlabel metal1 11500 12070 11500 12070 0 _046_
rlabel metal1 12834 10676 12834 10676 0 _047_
rlabel metal1 12144 10778 12144 10778 0 _048_
rlabel metal2 11086 7650 11086 7650 0 _049_
rlabel metal1 12006 9418 12006 9418 0 _050_
rlabel metal2 12328 10030 12328 10030 0 _051_
rlabel metal1 11914 10166 11914 10166 0 _052_
rlabel metal1 11684 11866 11684 11866 0 _053_
rlabel metal3 9522 12580 9522 12580 0 _054_
rlabel via2 4370 12699 4370 12699 0 _055_
rlabel metal1 4692 6290 4692 6290 0 _056_
rlabel metal1 5014 5134 5014 5134 0 _057_
rlabel metal2 5290 5576 5290 5576 0 _058_
rlabel metal1 5060 5542 5060 5542 0 _059_
rlabel metal1 5461 5338 5461 5338 0 _060_
rlabel metal2 5198 4828 5198 4828 0 _061_
rlabel metal1 5221 5270 5221 5270 0 _062_
rlabel metal1 6348 2958 6348 2958 0 _063_
rlabel metal1 5934 4114 5934 4114 0 _064_
rlabel metal1 6026 3978 6026 3978 0 _065_
rlabel metal1 6026 3604 6026 3604 0 _066_
rlabel metal1 5750 3162 5750 3162 0 _067_
rlabel metal2 5382 3876 5382 3876 0 _068_
rlabel metal1 5566 3468 5566 3468 0 _069_
rlabel metal1 5589 4114 5589 4114 0 _070_
rlabel metal2 4600 12716 4600 12716 0 _071_
rlabel metal2 4140 12716 4140 12716 0 _072_
rlabel metal1 3588 13226 3588 13226 0 _073_
rlabel metal2 4278 12988 4278 12988 0 _074_
rlabel metal2 5428 8228 5428 8228 0 _075_
rlabel metal1 4968 4046 4968 4046 0 _076_
rlabel metal1 5106 4624 5106 4624 0 _077_
rlabel metal2 5290 4012 5290 4012 0 _078_
rlabel metal1 4968 3706 4968 3706 0 _079_
rlabel metal1 4140 4046 4140 4046 0 _080_
rlabel metal1 11040 7446 11040 7446 0 _081_
rlabel metal1 10534 5814 10534 5814 0 _082_
rlabel metal2 11546 5610 11546 5610 0 _083_
rlabel via1 8502 6698 8502 6698 0 _084_
rlabel metal1 11408 4726 11408 4726 0 _085_
rlabel metal1 8694 4998 8694 4998 0 _086_
rlabel metal1 9032 5270 9032 5270 0 _087_
rlabel metal2 8326 7378 8326 7378 0 _088_
rlabel metal2 8970 5984 8970 5984 0 _089_
rlabel metal1 8326 7990 8326 7990 0 _090_
rlabel metal1 8372 8058 8372 8058 0 _091_
rlabel metal1 5152 6766 5152 6766 0 _092_
rlabel metal2 5382 7072 5382 7072 0 _093_
rlabel metal1 4232 7242 4232 7242 0 _094_
rlabel metal2 4278 7480 4278 7480 0 _095_
rlabel metal1 1564 9622 1564 9622 0 _096_
rlabel metal1 2484 9350 2484 9350 0 _097_
rlabel metal2 3358 9622 3358 9622 0 _098_
rlabel metal1 2369 9554 2369 9554 0 _099_
rlabel metal1 2392 6766 2392 6766 0 _100_
rlabel metal2 2254 8432 2254 8432 0 _101_
rlabel metal2 2898 5950 2898 5950 0 _102_
rlabel metal2 2530 6256 2530 6256 0 _103_
rlabel metal1 3772 5542 3772 5542 0 _104_
rlabel metal2 3358 5168 3358 5168 0 _105_
rlabel metal1 8924 4046 8924 4046 0 _106_
rlabel metal2 8142 4182 8142 4182 0 _107_
rlabel metal2 8786 3808 8786 3808 0 _108_
rlabel metal1 10350 4148 10350 4148 0 _109_
rlabel metal1 6716 5746 6716 5746 0 _110_
rlabel metal1 6854 5610 6854 5610 0 _111_
rlabel metal2 6670 5236 6670 5236 0 _112_
rlabel metal2 6578 6086 6578 6086 0 _113_
rlabel metal2 6854 7990 6854 7990 0 _114_
rlabel metal2 5566 9724 5566 9724 0 _115_
rlabel metal1 4876 9690 4876 9690 0 _116_
rlabel metal2 5934 9792 5934 9792 0 _117_
rlabel via1 6670 10234 6670 10234 0 _118_
rlabel metal1 6900 10030 6900 10030 0 _119_
rlabel metal2 7222 9792 7222 9792 0 _120_
rlabel metal2 8050 10370 8050 10370 0 _121_
rlabel metal1 8740 10710 8740 10710 0 _122_
rlabel metal2 9062 11356 9062 11356 0 _123_
rlabel metal2 8970 11084 8970 11084 0 _124_
rlabel metal1 9430 10642 9430 10642 0 _125_
rlabel metal1 9660 9554 9660 9554 0 _126_
rlabel metal2 9706 9860 9706 9860 0 _127_
rlabel metal1 8878 10438 8878 10438 0 _128_
rlabel metal1 9660 8942 9660 8942 0 _129_
rlabel metal1 9108 9690 9108 9690 0 _130_
rlabel metal2 9430 9860 9430 9860 0 _131_
rlabel metal1 8786 10540 8786 10540 0 _132_
rlabel metal1 8326 10608 8326 10608 0 _133_
rlabel metal2 7314 10234 7314 10234 0 _134_
rlabel metal1 6578 10064 6578 10064 0 _135_
rlabel metal1 6394 9588 6394 9588 0 _136_
rlabel metal1 6072 9418 6072 9418 0 _137_
rlabel metal2 6302 9146 6302 9146 0 _138_
rlabel metal1 7268 5882 7268 5882 0 _139_
rlabel metal1 9936 10234 9936 10234 0 _140_
rlabel metal2 8786 9792 8786 9792 0 _141_
rlabel metal1 6578 8976 6578 8976 0 _142_
rlabel metal1 6026 9588 6026 9588 0 _143_
rlabel metal2 6670 9214 6670 9214 0 _144_
rlabel metal1 11178 9146 11178 9146 0 _145_
rlabel metal1 10810 9588 10810 9588 0 _146_
rlabel metal1 8786 9894 8786 9894 0 _147_
rlabel metal2 9338 11883 9338 11883 0 _148_
rlabel metal2 9522 11866 9522 11866 0 _149_
rlabel metal1 7958 12240 7958 12240 0 _150_
rlabel metal2 7958 11900 7958 11900 0 _151_
rlabel metal1 5980 10710 5980 10710 0 _152_
rlabel metal1 4968 13226 4968 13226 0 _153_
rlabel metal1 5382 10030 5382 10030 0 _154_
rlabel metal2 4738 6596 4738 6596 0 _155_
rlabel metal1 6440 4454 6440 4454 0 _156_
rlabel metal2 7038 5950 7038 5950 0 _157_
rlabel metal2 6026 5882 6026 5882 0 _158_
rlabel metal2 12098 9826 12098 9826 0 _159_
rlabel metal2 10074 13022 10074 13022 0 _160_
rlabel metal2 9982 13158 9982 13158 0 _161_
rlabel metal1 6946 12784 6946 12784 0 _162_
rlabel metal2 7038 13090 7038 13090 0 _163_
rlabel metal1 6026 11662 6026 11662 0 _164_
rlabel metal1 5658 12682 5658 12682 0 _165_
rlabel metal2 5198 12517 5198 12517 0 _166_
rlabel metal1 4416 13362 4416 13362 0 _167_
rlabel metal1 6118 12410 6118 12410 0 _168_
rlabel metal2 4094 11679 4094 11679 0 _169_
rlabel metal2 4186 11934 4186 11934 0 _170_
rlabel metal1 3588 11662 3588 11662 0 _171_
rlabel metal1 5980 11730 5980 11730 0 _172_
rlabel metal3 5382 12580 5382 12580 0 _173_
rlabel metal1 4968 11050 4968 11050 0 _174_
rlabel metal1 4600 11322 4600 11322 0 _175_
rlabel metal2 6486 8177 6486 8177 0 clk
rlabel metal1 7544 6970 7544 6970 0 clknet_0_clk
rlabel metal2 1886 5746 1886 5746 0 clknet_1_0__leaf_clk
rlabel metal1 7728 2482 7728 2482 0 clknet_1_1__leaf_clk
rlabel metal1 11638 8942 11638 8942 0 counter\[0\]
rlabel metal1 1610 10574 1610 10574 0 counter\[10\]
rlabel metal1 3266 11798 3266 11798 0 counter\[11\]
rlabel metal1 1932 6698 1932 6698 0 counter\[12\]
rlabel metal1 6440 4998 6440 4998 0 counter\[13\]
rlabel metal1 8326 4522 8326 4522 0 counter\[14\]
rlabel metal1 10212 4114 10212 4114 0 counter\[15\]
rlabel metal1 12696 6970 12696 6970 0 counter\[1\]
rlabel metal2 12558 11220 12558 11220 0 counter\[2\]
rlabel metal2 11730 5236 11730 5236 0 counter\[3\]
rlabel metal2 9338 4828 9338 4828 0 counter\[4\]
rlabel metal1 8832 12818 8832 12818 0 counter\[5\]
rlabel metal1 8050 12750 8050 12750 0 counter\[6\]
rlabel metal1 7590 8058 7590 8058 0 counter\[7\]
rlabel viali 5395 11730 5395 11730 0 counter\[8\]
rlabel metal1 5428 10642 5428 10642 0 counter\[9\]
rlabel via1 12558 10098 12558 10098 0 net1
rlabel metal2 10350 9996 10350 9996 0 net10
rlabel metal1 8418 13464 8418 13464 0 net11
rlabel metal1 9568 13294 9568 13294 0 net12
rlabel metal1 8970 13838 8970 13838 0 net13
rlabel metal2 7222 13124 7222 13124 0 net14
rlabel metal1 9522 13770 9522 13770 0 net15
rlabel metal1 6716 13498 6716 13498 0 net16
rlabel metal2 12650 6834 12650 6834 0 net17
rlabel metal1 7866 2618 7866 2618 0 net18
rlabel metal1 2622 5610 2622 5610 0 net19
rlabel metal1 6072 13770 6072 13770 0 net2
rlabel metal2 10442 6800 10442 6800 0 net20
rlabel metal2 12742 8160 12742 8160 0 net21
rlabel metal2 8602 4590 8602 4590 0 net22
rlabel metal1 5474 6834 5474 6834 0 net23
rlabel metal1 5520 12614 5520 12614 0 net24
rlabel metal1 4692 3570 4692 3570 0 net25
rlabel metal1 2346 4522 2346 4522 0 net26
rlabel metal2 12006 6188 12006 6188 0 net27
rlabel metal1 11178 10030 11178 10030 0 net28
rlabel metal1 11707 10030 11707 10030 0 net29
rlabel metal1 5106 12750 5106 12750 0 net3
rlabel metal1 2438 6664 2438 6664 0 net4
rlabel metal1 5382 6222 5382 6222 0 net5
rlabel metal1 5842 2414 5842 2414 0 net6
rlabel metal1 6072 2890 6072 2890 0 net7
rlabel metal2 12466 10812 12466 10812 0 net8
rlabel metal1 12558 10030 12558 10030 0 net9
rlabel metal1 7222 2822 7222 2822 0 out
rlabel metal2 13018 9265 13018 9265 0 psc[0]
rlabel metal2 5290 14399 5290 14399 0 psc[10]
rlabel metal1 5980 13906 5980 13906 0 psc[11]
rlabel metal3 751 6188 751 6188 0 psc[12]
rlabel metal2 5198 1027 5198 1027 0 psc[13]
rlabel metal2 5842 1622 5842 1622 0 psc[14]
rlabel metal1 6624 3026 6624 3026 0 psc[15]
rlabel metal2 12926 10693 12926 10693 0 psc[1]
rlabel via2 12742 8925 12742 8925 0 psc[2]
rlabel metal2 12834 11033 12834 11033 0 psc[3]
rlabel metal1 9798 13906 9798 13906 0 psc[4]
rlabel metal1 9246 13906 9246 13906 0 psc[5]
rlabel metal1 7866 13906 7866 13906 0 psc[6]
rlabel metal1 7176 13906 7176 13906 0 psc[7]
rlabel metal1 8740 13974 8740 13974 0 psc[8]
rlabel metal1 6532 13906 6532 13906 0 psc[9]
rlabel via2 13018 3485 13018 3485 0 rst
<< properties >>
string FIXED_BBOX 0 0 14478 16622
<< end >>
