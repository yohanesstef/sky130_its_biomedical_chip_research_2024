magic
tech sky130A
magscale 1 2
timestamp 1730019635
<< error_p >>
rect -29 171 29 177
rect -29 137 -17 171
rect -29 131 29 137
<< nwell >>
rect -109 -224 109 190
<< pmos >>
rect -15 -162 15 90
<< pdiff >>
rect -73 78 -15 90
rect -73 -150 -61 78
rect -27 -150 -15 78
rect -73 -162 -15 -150
rect 15 78 73 90
rect 15 -150 27 78
rect 61 -150 73 78
rect 15 -162 73 -150
<< pdiffc >>
rect -61 -150 -27 78
rect 27 -150 61 78
<< poly >>
rect -33 171 33 187
rect -33 137 -17 171
rect 17 137 33 171
rect -33 121 33 137
rect -15 90 15 121
rect -15 -188 15 -162
<< polycont >>
rect -17 137 17 171
<< locali >>
rect -33 137 -17 171
rect 17 137 33 171
rect -61 78 -27 94
rect -61 -166 -27 -150
rect 27 78 61 94
rect 27 -166 61 -150
<< viali >>
rect -17 137 17 171
rect -61 -150 -27 78
rect 27 -150 61 78
<< metal1 >>
rect -29 171 29 177
rect -29 137 -17 171
rect 17 137 29 171
rect -29 131 29 137
rect -67 78 -21 90
rect -67 -150 -61 78
rect -27 -150 -21 78
rect -67 -162 -21 -150
rect 21 78 67 90
rect 21 -150 27 78
rect 61 -150 67 78
rect 21 -162 67 -150
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
