module freq_psc (clk,
    out,
    rst,
    psc);
 input clk;
 output out;
 input rst;
 input [31:0] psc;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire \psc_cnt[0] ;
 wire \psc_cnt[10] ;
 wire \psc_cnt[11] ;
 wire \psc_cnt[12] ;
 wire \psc_cnt[13] ;
 wire \psc_cnt[14] ;
 wire \psc_cnt[15] ;
 wire \psc_cnt[16] ;
 wire \psc_cnt[17] ;
 wire \psc_cnt[18] ;
 wire \psc_cnt[19] ;
 wire \psc_cnt[1] ;
 wire \psc_cnt[20] ;
 wire \psc_cnt[21] ;
 wire \psc_cnt[22] ;
 wire \psc_cnt[23] ;
 wire \psc_cnt[24] ;
 wire \psc_cnt[25] ;
 wire \psc_cnt[26] ;
 wire \psc_cnt[27] ;
 wire \psc_cnt[28] ;
 wire \psc_cnt[29] ;
 wire \psc_cnt[2] ;
 wire \psc_cnt[30] ;
 wire \psc_cnt[31] ;
 wire \psc_cnt[3] ;
 wire \psc_cnt[4] ;
 wire \psc_cnt[5] ;
 wire \psc_cnt[6] ;
 wire \psc_cnt[7] ;
 wire \psc_cnt[8] ;
 wire \psc_cnt[9] ;

 sky130_fd_sc_hd__inv_2 _236_ (.A(\psc_cnt[24] ),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _237_ (.A(psc[22]),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _238_ (.A(psc[21]),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _239_ (.A(\psc_cnt[20] ),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _240_ (.A(\psc_cnt[19] ),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _241_ (.A(psc[18]),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _242_ (.A(psc[17]),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _243_ (.A(psc[16]),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _244_ (.A(\psc_cnt[15] ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _245_ (.A(\psc_cnt[14] ),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _246_ (.A(\psc_cnt[13] ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _247_ (.A(\psc_cnt[12] ),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _248_ (.A(\psc_cnt[11] ),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _249_ (.A(\psc_cnt[10] ),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _250_ (.A(\psc_cnt[9] ),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _251_ (.A(\psc_cnt[8] ),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _252_ (.A(psc[8]),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _253_ (.A(psc[7]),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _254_ (.A(psc[6]),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _255_ (.A(psc[5]),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _256_ (.A(psc[4]),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _257_ (.A(psc[3]),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _258_ (.A(psc[2]),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _259_ (.A(psc[1]),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _260_ (.A(psc[0]),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _261_ (.A(\psc_cnt[25] ),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _262_ (.A(\psc_cnt[26] ),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _263_ (.A(\psc_cnt[28] ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _264_ (.A(\psc_cnt[29] ),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _265_ (.A(\psc_cnt[31] ),
    .Y(_095_));
 sky130_fd_sc_hd__inv_2 _266_ (.A(rst),
    .Y(_032_));
 sky130_fd_sc_hd__and2_2 _267_ (.A(psc[15]),
    .B(_074_),
    .X(_096_));
 sky130_fd_sc_hd__o22a_2 _268_ (.A1(psc[15]),
    .A2(_074_),
    .B1(psc[14]),
    .B2(_075_),
    .X(_097_));
 sky130_fd_sc_hd__a22oi_2 _269_ (.A1(psc[14]),
    .A2(_075_),
    .B1(psc[13]),
    .B2(_076_),
    .Y(_098_));
 sky130_fd_sc_hd__o22a_2 _270_ (.A1(psc[13]),
    .A2(_076_),
    .B1(_077_),
    .B2(psc[12]),
    .X(_099_));
 sky130_fd_sc_hd__nand2b_2 _271_ (.A_N(_099_),
    .B(_098_),
    .Y(_100_));
 sky130_fd_sc_hd__a21oi_2 _272_ (.A1(_097_),
    .A2(_100_),
    .B1(_096_),
    .Y(_101_));
 sky130_fd_sc_hd__a21oi_2 _273_ (.A1(_077_),
    .A2(psc[12]),
    .B1(_096_),
    .Y(_102_));
 sky130_fd_sc_hd__and4_2 _274_ (.A(_097_),
    .B(_098_),
    .C(_099_),
    .D(_102_),
    .X(_103_));
 sky130_fd_sc_hd__and2b_2 _275_ (.A_N(\psc_cnt[11] ),
    .B(psc[11]),
    .X(_104_));
 sky130_fd_sc_hd__o22a_2 _276_ (.A1(psc[11]),
    .A2(_078_),
    .B1(psc[10]),
    .B2(_079_),
    .X(_105_));
 sky130_fd_sc_hd__a221oi_2 _277_ (.A1(psc[10]),
    .A2(_079_),
    .B1(psc[9]),
    .B2(_080_),
    .C1(_104_),
    .Y(_106_));
 sky130_fd_sc_hd__nand2_2 _278_ (.A(_105_),
    .B(_106_),
    .Y(_107_));
 sky130_fd_sc_hd__o22a_2 _279_ (.A1(psc[9]),
    .A2(_080_),
    .B1(_081_),
    .B2(psc[8]),
    .X(_108_));
 sky130_fd_sc_hd__a22o_2 _280_ (.A1(_085_),
    .A2(\psc_cnt[5] ),
    .B1(\psc_cnt[4] ),
    .B2(_086_),
    .X(_109_));
 sky130_fd_sc_hd__a211o_2 _281_ (.A1(_089_),
    .A2(\psc_cnt[1] ),
    .B1(_090_),
    .C1(\psc_cnt[0] ),
    .X(_110_));
 sky130_fd_sc_hd__o22a_2 _282_ (.A1(_088_),
    .A2(\psc_cnt[2] ),
    .B1(_089_),
    .B2(\psc_cnt[1] ),
    .X(_111_));
 sky130_fd_sc_hd__a22o_2 _283_ (.A1(_087_),
    .A2(\psc_cnt[3] ),
    .B1(_088_),
    .B2(\psc_cnt[2] ),
    .X(_112_));
 sky130_fd_sc_hd__a21o_2 _284_ (.A1(_110_),
    .A2(_111_),
    .B1(_112_),
    .X(_113_));
 sky130_fd_sc_hd__o22a_2 _285_ (.A1(\psc_cnt[4] ),
    .A2(_086_),
    .B1(_087_),
    .B2(\psc_cnt[3] ),
    .X(_114_));
 sky130_fd_sc_hd__a21o_2 _286_ (.A1(_113_),
    .A2(_114_),
    .B1(_109_),
    .X(_115_));
 sky130_fd_sc_hd__o22a_2 _287_ (.A1(_084_),
    .A2(\psc_cnt[6] ),
    .B1(_085_),
    .B2(\psc_cnt[5] ),
    .X(_116_));
 sky130_fd_sc_hd__a22o_2 _288_ (.A1(_083_),
    .A2(\psc_cnt[7] ),
    .B1(_084_),
    .B2(\psc_cnt[6] ),
    .X(_117_));
 sky130_fd_sc_hd__a21o_2 _289_ (.A1(_115_),
    .A2(_116_),
    .B1(_117_),
    .X(_118_));
 sky130_fd_sc_hd__o221a_2 _290_ (.A1(\psc_cnt[8] ),
    .A2(_082_),
    .B1(_083_),
    .B2(\psc_cnt[7] ),
    .C1(_108_),
    .X(_119_));
 sky130_fd_sc_hd__and4_2 _291_ (.A(_103_),
    .B(_105_),
    .C(_106_),
    .D(_119_),
    .X(_120_));
 sky130_fd_sc_hd__o22a_2 _292_ (.A1(_104_),
    .A2(_105_),
    .B1(_107_),
    .B2(_108_),
    .X(_121_));
 sky130_fd_sc_hd__and2b_2 _293_ (.A_N(_121_),
    .B(_103_),
    .X(_122_));
 sky130_fd_sc_hd__a211o_2 _294_ (.A1(_118_),
    .A2(_120_),
    .B1(_122_),
    .C1(_101_),
    .X(_123_));
 sky130_fd_sc_hd__a2bb2o_2 _295_ (.A1_N(psc[19]),
    .A2_N(_070_),
    .B1(_071_),
    .B2(\psc_cnt[18] ),
    .X(_124_));
 sky130_fd_sc_hd__nand2_2 _296_ (.A(psc[19]),
    .B(_070_),
    .Y(_125_));
 sky130_fd_sc_hd__or2_2 _297_ (.A(_071_),
    .B(\psc_cnt[18] ),
    .X(_126_));
 sky130_fd_sc_hd__and3b_2 _298_ (.A_N(_124_),
    .B(_125_),
    .C(_126_),
    .X(_127_));
 sky130_fd_sc_hd__a22o_2 _299_ (.A1(_072_),
    .A2(\psc_cnt[17] ),
    .B1(\psc_cnt[16] ),
    .B2(_073_),
    .X(_128_));
 sky130_fd_sc_hd__or2_2 _300_ (.A(_072_),
    .B(\psc_cnt[17] ),
    .X(_129_));
 sky130_fd_sc_hd__o21a_2 _301_ (.A1(\psc_cnt[16] ),
    .A2(_073_),
    .B1(_127_),
    .X(_130_));
 sky130_fd_sc_hd__and2b_2 _302_ (.A_N(psc[23]),
    .B(\psc_cnt[23] ),
    .X(_131_));
 sky130_fd_sc_hd__a21o_2 _303_ (.A1(_067_),
    .A2(\psc_cnt[22] ),
    .B1(_131_),
    .X(_132_));
 sky130_fd_sc_hd__and2b_2 _304_ (.A_N(psc[20]),
    .B(\psc_cnt[20] ),
    .X(_133_));
 sky130_fd_sc_hd__and2b_2 _305_ (.A_N(psc[21]),
    .B(\psc_cnt[21] ),
    .X(_134_));
 sky130_fd_sc_hd__a2111o_2 _306_ (.A1(_067_),
    .A2(\psc_cnt[22] ),
    .B1(_131_),
    .C1(_133_),
    .D1(_134_),
    .X(_135_));
 sky130_fd_sc_hd__and2b_2 _307_ (.A_N(psc[27]),
    .B(\psc_cnt[27] ),
    .X(_136_));
 sky130_fd_sc_hd__and2b_2 _308_ (.A_N(psc[26]),
    .B(\psc_cnt[26] ),
    .X(_137_));
 sky130_fd_sc_hd__nor2_2 _309_ (.A(_136_),
    .B(_137_),
    .Y(_138_));
 sky130_fd_sc_hd__and2b_2 _310_ (.A_N(\psc_cnt[27] ),
    .B(psc[27]),
    .X(_139_));
 sky130_fd_sc_hd__and2b_2 _311_ (.A_N(\psc_cnt[26] ),
    .B(psc[26]),
    .X(_140_));
 sky130_fd_sc_hd__or4_2 _312_ (.A(_136_),
    .B(_137_),
    .C(_139_),
    .D(_140_),
    .X(_141_));
 sky130_fd_sc_hd__and2b_2 _313_ (.A_N(\psc_cnt[24] ),
    .B(psc[24]),
    .X(_142_));
 sky130_fd_sc_hd__and2b_2 _314_ (.A_N(\psc_cnt[25] ),
    .B(psc[25]),
    .X(_143_));
 sky130_fd_sc_hd__and2b_2 _315_ (.A_N(\psc_cnt[23] ),
    .B(psc[23]),
    .X(_144_));
 sky130_fd_sc_hd__or3_2 _316_ (.A(_142_),
    .B(_143_),
    .C(_144_),
    .X(_145_));
 sky130_fd_sc_hd__or3_2 _317_ (.A(_135_),
    .B(_141_),
    .C(_145_),
    .X(_146_));
 sky130_fd_sc_hd__and2b_2 _318_ (.A_N(psc[31]),
    .B(\psc_cnt[31] ),
    .X(_147_));
 sky130_fd_sc_hd__and2b_2 _319_ (.A_N(psc[30]),
    .B(\psc_cnt[30] ),
    .X(_148_));
 sky130_fd_sc_hd__nor2_2 _320_ (.A(_147_),
    .B(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__and2b_2 _321_ (.A_N(\psc_cnt[31] ),
    .B(psc[31]),
    .X(_150_));
 sky130_fd_sc_hd__and2b_2 _322_ (.A_N(\psc_cnt[30] ),
    .B(psc[30]),
    .X(_151_));
 sky130_fd_sc_hd__and2_2 _323_ (.A(_094_),
    .B(psc[29]),
    .X(_152_));
 sky130_fd_sc_hd__or4_2 _324_ (.A(_147_),
    .B(_148_),
    .C(_150_),
    .D(_151_),
    .X(_153_));
 sky130_fd_sc_hd__nor2_2 _325_ (.A(_152_),
    .B(_153_),
    .Y(_154_));
 sky130_fd_sc_hd__o22a_2 _326_ (.A1(_094_),
    .A2(psc[29]),
    .B1(psc[28]),
    .B2(_093_),
    .X(_155_));
 sky130_fd_sc_hd__and2b_2 _327_ (.A_N(\psc_cnt[28] ),
    .B(psc[28]),
    .X(_156_));
 sky130_fd_sc_hd__a21oi_2 _328_ (.A1(_069_),
    .A2(psc[20]),
    .B1(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__o22a_2 _329_ (.A1(_066_),
    .A2(psc[24]),
    .B1(_091_),
    .B2(psc[25]),
    .X(_158_));
 sky130_fd_sc_hd__o22a_2 _330_ (.A1(_067_),
    .A2(\psc_cnt[22] ),
    .B1(_068_),
    .B2(\psc_cnt[21] ),
    .X(_159_));
 sky130_fd_sc_hd__and4_2 _331_ (.A(_155_),
    .B(_157_),
    .C(_158_),
    .D(_159_),
    .X(_160_));
 sky130_fd_sc_hd__or4b_2 _332_ (.A(_152_),
    .B(_153_),
    .C(_156_),
    .D_N(_155_),
    .X(_161_));
 sky130_fd_sc_hd__or4_2 _333_ (.A(_141_),
    .B(_142_),
    .C(_143_),
    .D(_161_),
    .X(_162_));
 sky130_fd_sc_hd__and3b_2 _334_ (.A_N(_146_),
    .B(_154_),
    .C(_160_),
    .X(_163_));
 sky130_fd_sc_hd__and4b_2 _335_ (.A_N(_128_),
    .B(_129_),
    .C(_130_),
    .D(_163_),
    .X(_164_));
 sky130_fd_sc_hd__a32o_2 _336_ (.A1(_127_),
    .A2(_128_),
    .A3(_129_),
    .B1(_125_),
    .B2(_124_),
    .X(_165_));
 sky130_fd_sc_hd__and2_2 _337_ (.A(_163_),
    .B(_165_),
    .X(_166_));
 sky130_fd_sc_hd__o32a_2 _338_ (.A1(_141_),
    .A2(_143_),
    .A3(_158_),
    .B1(_139_),
    .B2(_138_),
    .X(_167_));
 sky130_fd_sc_hd__o32a_2 _339_ (.A1(_152_),
    .A2(_153_),
    .A3(_155_),
    .B1(_150_),
    .B2(_149_),
    .X(_168_));
 sky130_fd_sc_hd__o21ai_2 _340_ (.A1(_161_),
    .A2(_167_),
    .B1(_168_),
    .Y(_169_));
 sky130_fd_sc_hd__o21ba_2 _341_ (.A1(_132_),
    .A2(_159_),
    .B1_N(_144_),
    .X(_170_));
 sky130_fd_sc_hd__and4b_2 _342_ (.A_N(_162_),
    .B(_135_),
    .C(_158_),
    .D(_170_),
    .X(_171_));
 sky130_fd_sc_hd__or3_2 _343_ (.A(_166_),
    .B(_169_),
    .C(_171_),
    .X(_172_));
 sky130_fd_sc_hd__a21oi_2 _344_ (.A1(_123_),
    .A2(_164_),
    .B1(_172_),
    .Y(_173_));
 sky130_fd_sc_hd__xnor2_2 _345_ (.A(out),
    .B(_173_),
    .Y(_065_));
 sky130_fd_sc_hd__and2b_2 _346_ (.A_N(\psc_cnt[0] ),
    .B(_173_),
    .X(_000_));
 sky130_fd_sc_hd__or2_2 _347_ (.A(\psc_cnt[1] ),
    .B(\psc_cnt[0] ),
    .X(_174_));
 sky130_fd_sc_hd__nand2_2 _348_ (.A(\psc_cnt[1] ),
    .B(\psc_cnt[0] ),
    .Y(_175_));
 sky130_fd_sc_hd__and3_2 _349_ (.A(_173_),
    .B(_174_),
    .C(_175_),
    .X(_011_));
 sky130_fd_sc_hd__a21o_2 _350_ (.A1(\psc_cnt[1] ),
    .A2(\psc_cnt[0] ),
    .B1(\psc_cnt[2] ),
    .X(_176_));
 sky130_fd_sc_hd__nand3_2 _351_ (.A(\psc_cnt[2] ),
    .B(\psc_cnt[1] ),
    .C(\psc_cnt[0] ),
    .Y(_177_));
 sky130_fd_sc_hd__and3_2 _352_ (.A(_173_),
    .B(_176_),
    .C(_177_),
    .X(_022_));
 sky130_fd_sc_hd__a31o_2 _353_ (.A1(\psc_cnt[2] ),
    .A2(\psc_cnt[1] ),
    .A3(\psc_cnt[0] ),
    .B1(\psc_cnt[3] ),
    .X(_178_));
 sky130_fd_sc_hd__and4_2 _354_ (.A(\psc_cnt[3] ),
    .B(\psc_cnt[2] ),
    .C(\psc_cnt[1] ),
    .D(\psc_cnt[0] ),
    .X(_179_));
 sky130_fd_sc_hd__and3b_2 _355_ (.A_N(_179_),
    .B(_173_),
    .C(_178_),
    .X(_025_));
 sky130_fd_sc_hd__or2_2 _356_ (.A(\psc_cnt[4] ),
    .B(_179_),
    .X(_180_));
 sky130_fd_sc_hd__nand2_2 _357_ (.A(\psc_cnt[4] ),
    .B(_179_),
    .Y(_181_));
 sky130_fd_sc_hd__and3_2 _358_ (.A(_173_),
    .B(_180_),
    .C(_181_),
    .X(_026_));
 sky130_fd_sc_hd__a21o_2 _359_ (.A1(\psc_cnt[4] ),
    .A2(_179_),
    .B1(\psc_cnt[5] ),
    .X(_182_));
 sky130_fd_sc_hd__and2_2 _360_ (.A(\psc_cnt[5] ),
    .B(\psc_cnt[4] ),
    .X(_183_));
 sky130_fd_sc_hd__and2_2 _361_ (.A(_179_),
    .B(_183_),
    .X(_184_));
 sky130_fd_sc_hd__and3b_2 _362_ (.A_N(_184_),
    .B(_173_),
    .C(_182_),
    .X(_027_));
 sky130_fd_sc_hd__or2_2 _363_ (.A(\psc_cnt[6] ),
    .B(_184_),
    .X(_185_));
 sky130_fd_sc_hd__nand2_2 _364_ (.A(\psc_cnt[6] ),
    .B(_184_),
    .Y(_186_));
 sky130_fd_sc_hd__and3_2 _365_ (.A(_173_),
    .B(_185_),
    .C(_186_),
    .X(_028_));
 sky130_fd_sc_hd__a31o_2 _366_ (.A1(\psc_cnt[6] ),
    .A2(_179_),
    .A3(_183_),
    .B1(\psc_cnt[7] ),
    .X(_187_));
 sky130_fd_sc_hd__and4_2 _367_ (.A(\psc_cnt[7] ),
    .B(\psc_cnt[6] ),
    .C(_179_),
    .D(_183_),
    .X(_188_));
 sky130_fd_sc_hd__and3b_2 _368_ (.A_N(_188_),
    .B(_173_),
    .C(_187_),
    .X(_029_));
 sky130_fd_sc_hd__or2_2 _369_ (.A(\psc_cnt[8] ),
    .B(_188_),
    .X(_189_));
 sky130_fd_sc_hd__nand2_2 _370_ (.A(\psc_cnt[8] ),
    .B(_188_),
    .Y(_190_));
 sky130_fd_sc_hd__and3_2 _371_ (.A(_173_),
    .B(_189_),
    .C(_190_),
    .X(_030_));
 sky130_fd_sc_hd__nand2_2 _372_ (.A(_080_),
    .B(_190_),
    .Y(_191_));
 sky130_fd_sc_hd__nor2_2 _373_ (.A(_080_),
    .B(_081_),
    .Y(_192_));
 sky130_fd_sc_hd__and2_2 _374_ (.A(_188_),
    .B(_192_),
    .X(_193_));
 sky130_fd_sc_hd__and3b_2 _375_ (.A_N(_193_),
    .B(_173_),
    .C(_191_),
    .X(_031_));
 sky130_fd_sc_hd__or2_2 _376_ (.A(\psc_cnt[10] ),
    .B(_193_),
    .X(_194_));
 sky130_fd_sc_hd__and3_2 _377_ (.A(\psc_cnt[10] ),
    .B(_188_),
    .C(_192_),
    .X(_195_));
 sky130_fd_sc_hd__and3b_2 _378_ (.A_N(_195_),
    .B(_173_),
    .C(_194_),
    .X(_001_));
 sky130_fd_sc_hd__or2_2 _379_ (.A(\psc_cnt[11] ),
    .B(_195_),
    .X(_196_));
 sky130_fd_sc_hd__and4_2 _380_ (.A(\psc_cnt[11] ),
    .B(\psc_cnt[10] ),
    .C(_188_),
    .D(_192_),
    .X(_197_));
 sky130_fd_sc_hd__and3b_2 _381_ (.A_N(_197_),
    .B(_173_),
    .C(_196_),
    .X(_002_));
 sky130_fd_sc_hd__and2_2 _382_ (.A(\psc_cnt[12] ),
    .B(_197_),
    .X(_198_));
 sky130_fd_sc_hd__or2_2 _383_ (.A(\psc_cnt[12] ),
    .B(_197_),
    .X(_199_));
 sky130_fd_sc_hd__and3b_2 _384_ (.A_N(_198_),
    .B(_199_),
    .C(_173_),
    .X(_003_));
 sky130_fd_sc_hd__or2_2 _385_ (.A(\psc_cnt[13] ),
    .B(_198_),
    .X(_200_));
 sky130_fd_sc_hd__and3_2 _386_ (.A(\psc_cnt[13] ),
    .B(\psc_cnt[12] ),
    .C(_197_),
    .X(_201_));
 sky130_fd_sc_hd__and3b_2 _387_ (.A_N(_201_),
    .B(_173_),
    .C(_200_),
    .X(_004_));
 sky130_fd_sc_hd__or2_2 _388_ (.A(\psc_cnt[14] ),
    .B(_201_),
    .X(_202_));
 sky130_fd_sc_hd__nand2_2 _389_ (.A(\psc_cnt[14] ),
    .B(_201_),
    .Y(_203_));
 sky130_fd_sc_hd__and3_2 _390_ (.A(_173_),
    .B(_202_),
    .C(_203_),
    .X(_005_));
 sky130_fd_sc_hd__nor2_2 _391_ (.A(_074_),
    .B(_075_),
    .Y(_204_));
 sky130_fd_sc_hd__and4_2 _392_ (.A(\psc_cnt[13] ),
    .B(\psc_cnt[12] ),
    .C(_197_),
    .D(_204_),
    .X(_205_));
 sky130_fd_sc_hd__nand2_2 _393_ (.A(_074_),
    .B(_203_),
    .Y(_206_));
 sky130_fd_sc_hd__and3b_2 _394_ (.A_N(_205_),
    .B(_206_),
    .C(_173_),
    .X(_006_));
 sky130_fd_sc_hd__or2_2 _395_ (.A(\psc_cnt[16] ),
    .B(_205_),
    .X(_207_));
 sky130_fd_sc_hd__and2_2 _396_ (.A(\psc_cnt[16] ),
    .B(_205_),
    .X(_208_));
 sky130_fd_sc_hd__and3b_2 _397_ (.A_N(_208_),
    .B(_173_),
    .C(_207_),
    .X(_007_));
 sky130_fd_sc_hd__and3_2 _398_ (.A(\psc_cnt[17] ),
    .B(\psc_cnt[16] ),
    .C(_205_),
    .X(_209_));
 sky130_fd_sc_hd__or2_2 _399_ (.A(\psc_cnt[17] ),
    .B(_208_),
    .X(_210_));
 sky130_fd_sc_hd__and3b_2 _400_ (.A_N(_209_),
    .B(_210_),
    .C(_173_),
    .X(_008_));
 sky130_fd_sc_hd__nand2_2 _401_ (.A(\psc_cnt[18] ),
    .B(_209_),
    .Y(_211_));
 sky130_fd_sc_hd__o211a_2 _402_ (.A1(\psc_cnt[18] ),
    .A2(_209_),
    .B1(_211_),
    .C1(_173_),
    .X(_009_));
 sky130_fd_sc_hd__nand2_2 _403_ (.A(_070_),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__and4_2 _404_ (.A(\psc_cnt[19] ),
    .B(\psc_cnt[18] ),
    .C(\psc_cnt[17] ),
    .D(\psc_cnt[16] ),
    .X(_213_));
 sky130_fd_sc_hd__and2_2 _405_ (.A(_205_),
    .B(_213_),
    .X(_214_));
 sky130_fd_sc_hd__and3b_2 _406_ (.A_N(_214_),
    .B(_173_),
    .C(_212_),
    .X(_010_));
 sky130_fd_sc_hd__or2_2 _407_ (.A(\psc_cnt[20] ),
    .B(_214_),
    .X(_215_));
 sky130_fd_sc_hd__and3_2 _408_ (.A(\psc_cnt[20] ),
    .B(_205_),
    .C(_213_),
    .X(_216_));
 sky130_fd_sc_hd__and3b_2 _409_ (.A_N(_216_),
    .B(_173_),
    .C(_215_),
    .X(_012_));
 sky130_fd_sc_hd__nand2_2 _410_ (.A(\psc_cnt[21] ),
    .B(_216_),
    .Y(_217_));
 sky130_fd_sc_hd__o211a_2 _411_ (.A1(\psc_cnt[21] ),
    .A2(_216_),
    .B1(_217_),
    .C1(_173_),
    .X(_013_));
 sky130_fd_sc_hd__a21o_2 _412_ (.A1(\psc_cnt[21] ),
    .A2(_216_),
    .B1(\psc_cnt[22] ),
    .X(_218_));
 sky130_fd_sc_hd__and3_2 _413_ (.A(\psc_cnt[22] ),
    .B(\psc_cnt[21] ),
    .C(\psc_cnt[20] ),
    .X(_219_));
 sky130_fd_sc_hd__nand2_2 _414_ (.A(_214_),
    .B(_219_),
    .Y(_220_));
 sky130_fd_sc_hd__and3_2 _415_ (.A(_173_),
    .B(_218_),
    .C(_220_),
    .X(_014_));
 sky130_fd_sc_hd__a31o_2 _416_ (.A1(_205_),
    .A2(_213_),
    .A3(_219_),
    .B1(\psc_cnt[23] ),
    .X(_221_));
 sky130_fd_sc_hd__and3_2 _417_ (.A(\psc_cnt[23] ),
    .B(_213_),
    .C(_219_),
    .X(_222_));
 sky130_fd_sc_hd__and2_2 _418_ (.A(_205_),
    .B(_222_),
    .X(_223_));
 sky130_fd_sc_hd__and3b_2 _419_ (.A_N(_223_),
    .B(_173_),
    .C(_221_),
    .X(_015_));
 sky130_fd_sc_hd__or2_2 _420_ (.A(\psc_cnt[24] ),
    .B(_223_),
    .X(_224_));
 sky130_fd_sc_hd__and3_2 _421_ (.A(\psc_cnt[24] ),
    .B(_205_),
    .C(_222_),
    .X(_225_));
 sky130_fd_sc_hd__and3b_2 _422_ (.A_N(_225_),
    .B(_173_),
    .C(_224_),
    .X(_016_));
 sky130_fd_sc_hd__nand2_2 _423_ (.A(\psc_cnt[25] ),
    .B(_225_),
    .Y(_226_));
 sky130_fd_sc_hd__o211a_2 _424_ (.A1(\psc_cnt[25] ),
    .A2(_225_),
    .B1(_226_),
    .C1(_173_),
    .X(_017_));
 sky130_fd_sc_hd__nand2_2 _425_ (.A(_092_),
    .B(_226_),
    .Y(_227_));
 sky130_fd_sc_hd__o211a_2 _426_ (.A1(_092_),
    .A2(_226_),
    .B1(_227_),
    .C1(_173_),
    .X(_018_));
 sky130_fd_sc_hd__a31o_2 _427_ (.A1(\psc_cnt[25] ),
    .A2(\psc_cnt[26] ),
    .A3(_225_),
    .B1(\psc_cnt[27] ),
    .X(_228_));
 sky130_fd_sc_hd__and4_2 _428_ (.A(\psc_cnt[24] ),
    .B(\psc_cnt[25] ),
    .C(\psc_cnt[26] ),
    .D(\psc_cnt[27] ),
    .X(_229_));
 sky130_fd_sc_hd__and3_2 _429_ (.A(_205_),
    .B(_222_),
    .C(_229_),
    .X(_230_));
 sky130_fd_sc_hd__and3b_2 _430_ (.A_N(_230_),
    .B(_173_),
    .C(_228_),
    .X(_019_));
 sky130_fd_sc_hd__nand2_2 _431_ (.A(\psc_cnt[28] ),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__o211a_2 _432_ (.A1(\psc_cnt[28] ),
    .A2(_230_),
    .B1(_231_),
    .C1(_173_),
    .X(_020_));
 sky130_fd_sc_hd__nand2_2 _433_ (.A(_094_),
    .B(_231_),
    .Y(_232_));
 sky130_fd_sc_hd__and3_2 _434_ (.A(\psc_cnt[28] ),
    .B(\psc_cnt[29] ),
    .C(_230_),
    .X(_233_));
 sky130_fd_sc_hd__and3b_2 _435_ (.A_N(_233_),
    .B(_173_),
    .C(_232_),
    .X(_021_));
 sky130_fd_sc_hd__or2_2 _436_ (.A(\psc_cnt[30] ),
    .B(_233_),
    .X(_234_));
 sky130_fd_sc_hd__nand2_2 _437_ (.A(\psc_cnt[30] ),
    .B(_233_),
    .Y(_235_));
 sky130_fd_sc_hd__and3_2 _438_ (.A(_173_),
    .B(_234_),
    .C(_235_),
    .X(_023_));
 sky130_fd_sc_hd__a21boi_2 _439_ (.A1(_095_),
    .A2(_235_),
    .B1_N(_173_),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _440_ (.A(rst),
    .Y(_033_));
 sky130_fd_sc_hd__inv_2 _441_ (.A(rst),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _442_ (.A(rst),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _443_ (.A(rst),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _444_ (.A(rst),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _445_ (.A(rst),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _446_ (.A(rst),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _447_ (.A(rst),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _448_ (.A(rst),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _449_ (.A(rst),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _450_ (.A(rst),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _451_ (.A(rst),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _452_ (.A(rst),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _453_ (.A(rst),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _454_ (.A(rst),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _455_ (.A(rst),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _456_ (.A(rst),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _457_ (.A(rst),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _458_ (.A(rst),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _459_ (.A(rst),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _460_ (.A(rst),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _461_ (.A(rst),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _462_ (.A(rst),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _463_ (.A(rst),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _464_ (.A(rst),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _465_ (.A(rst),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _466_ (.A(rst),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _467_ (.A(rst),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _468_ (.A(rst),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _469_ (.A(rst),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _470_ (.A(rst),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _471_ (.A(rst),
    .Y(_064_));
 sky130_fd_sc_hd__dfrtp_2 _472_ (.CLK(clk),
    .D(_000_),
    .RESET_B(_032_),
    .Q(\psc_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _473_ (.CLK(clk),
    .D(_011_),
    .RESET_B(_033_),
    .Q(\psc_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_2 _474_ (.CLK(clk),
    .D(_022_),
    .RESET_B(_034_),
    .Q(\psc_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _475_ (.CLK(clk),
    .D(_025_),
    .RESET_B(_035_),
    .Q(\psc_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_2 _476_ (.CLK(clk),
    .D(_026_),
    .RESET_B(_036_),
    .Q(\psc_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _477_ (.CLK(clk),
    .D(_027_),
    .RESET_B(_037_),
    .Q(\psc_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _478_ (.CLK(clk),
    .D(_028_),
    .RESET_B(_038_),
    .Q(\psc_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_2 _479_ (.CLK(clk),
    .D(_029_),
    .RESET_B(_039_),
    .Q(\psc_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_2 _480_ (.CLK(clk),
    .D(_030_),
    .RESET_B(_040_),
    .Q(\psc_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_2 _481_ (.CLK(clk),
    .D(_031_),
    .RESET_B(_041_),
    .Q(\psc_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_2 _482_ (.CLK(clk),
    .D(_001_),
    .RESET_B(_042_),
    .Q(\psc_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_2 _483_ (.CLK(clk),
    .D(_002_),
    .RESET_B(_043_),
    .Q(\psc_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_2 _484_ (.CLK(clk),
    .D(_003_),
    .RESET_B(_044_),
    .Q(\psc_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_2 _485_ (.CLK(clk),
    .D(_004_),
    .RESET_B(_045_),
    .Q(\psc_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_2 _486_ (.CLK(clk),
    .D(_005_),
    .RESET_B(_046_),
    .Q(\psc_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_2 _487_ (.CLK(clk),
    .D(_006_),
    .RESET_B(_047_),
    .Q(\psc_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_2 _488_ (.CLK(clk),
    .D(_007_),
    .RESET_B(_048_),
    .Q(\psc_cnt[16] ));
 sky130_fd_sc_hd__dfrtp_2 _489_ (.CLK(clk),
    .D(_008_),
    .RESET_B(_049_),
    .Q(\psc_cnt[17] ));
 sky130_fd_sc_hd__dfrtp_2 _490_ (.CLK(clk),
    .D(_009_),
    .RESET_B(_050_),
    .Q(\psc_cnt[18] ));
 sky130_fd_sc_hd__dfrtp_2 _491_ (.CLK(clk),
    .D(_010_),
    .RESET_B(_051_),
    .Q(\psc_cnt[19] ));
 sky130_fd_sc_hd__dfrtp_2 _492_ (.CLK(clk),
    .D(_012_),
    .RESET_B(_052_),
    .Q(\psc_cnt[20] ));
 sky130_fd_sc_hd__dfrtp_2 _493_ (.CLK(clk),
    .D(_013_),
    .RESET_B(_053_),
    .Q(\psc_cnt[21] ));
 sky130_fd_sc_hd__dfrtp_2 _494_ (.CLK(clk),
    .D(_014_),
    .RESET_B(_054_),
    .Q(\psc_cnt[22] ));
 sky130_fd_sc_hd__dfrtp_2 _495_ (.CLK(clk),
    .D(_015_),
    .RESET_B(_055_),
    .Q(\psc_cnt[23] ));
 sky130_fd_sc_hd__dfrtp_2 _496_ (.CLK(clk),
    .D(_016_),
    .RESET_B(_056_),
    .Q(\psc_cnt[24] ));
 sky130_fd_sc_hd__dfrtp_2 _497_ (.CLK(clk),
    .D(_017_),
    .RESET_B(_057_),
    .Q(\psc_cnt[25] ));
 sky130_fd_sc_hd__dfrtp_2 _498_ (.CLK(clk),
    .D(_018_),
    .RESET_B(_058_),
    .Q(\psc_cnt[26] ));
 sky130_fd_sc_hd__dfrtp_2 _499_ (.CLK(clk),
    .D(_019_),
    .RESET_B(_059_),
    .Q(\psc_cnt[27] ));
 sky130_fd_sc_hd__dfrtp_2 _500_ (.CLK(clk),
    .D(_020_),
    .RESET_B(_060_),
    .Q(\psc_cnt[28] ));
 sky130_fd_sc_hd__dfrtp_2 _501_ (.CLK(clk),
    .D(_021_),
    .RESET_B(_061_),
    .Q(\psc_cnt[29] ));
 sky130_fd_sc_hd__dfrtp_2 _502_ (.CLK(clk),
    .D(_023_),
    .RESET_B(_062_),
    .Q(\psc_cnt[30] ));
 sky130_fd_sc_hd__dfrtp_2 _503_ (.CLK(clk),
    .D(_024_),
    .RESET_B(_063_),
    .Q(\psc_cnt[31] ));
 sky130_fd_sc_hd__dfrtp_2 _504_ (.CLK(clk),
    .D(_065_),
    .RESET_B(_064_),
    .Q(out));
endmodule
