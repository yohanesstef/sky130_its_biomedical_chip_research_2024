magic
tech sky130A
magscale 1 2
timestamp 1729851530
<< error_p >>
rect -32 -491 32 -485
rect -32 -525 -20 -491
rect -32 -531 32 -525
<< nwell >>
rect -130 -544 130 578
<< pmos >>
rect -36 -444 36 516
<< pdiff >>
rect -94 504 -36 516
rect -94 -432 -82 504
rect -48 -432 -36 504
rect -94 -444 -36 -432
rect 36 504 94 516
rect 36 -432 48 504
rect 82 -432 94 504
rect 36 -444 94 -432
<< pdiffc >>
rect -82 -432 -48 504
rect 48 -432 82 504
<< poly >>
rect -36 516 36 542
rect -36 -491 36 -444
rect -36 -525 -20 -491
rect 20 -525 36 -491
rect -36 -541 36 -525
<< polycont >>
rect -20 -525 20 -491
<< locali >>
rect -82 504 -48 520
rect -82 -448 -48 -432
rect 48 504 82 520
rect 48 -448 82 -432
rect -36 -525 -20 -491
rect 20 -525 36 -491
<< viali >>
rect -82 -432 -48 504
rect 48 -432 82 504
rect -20 -525 20 -491
<< metal1 >>
rect -88 504 -42 516
rect -88 -432 -82 504
rect -48 -432 -42 504
rect -88 -444 -42 -432
rect 42 504 88 516
rect 42 -432 48 504
rect 82 -432 88 504
rect 42 -444 88 -432
rect -32 -491 32 -485
rect -32 -525 -20 -491
rect 20 -525 32 -491
rect -32 -531 32 -525
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.8 l 0.36 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
