magic
tech sky130A
magscale 1 2
timestamp 1730527170
<< nwell >>
rect -943 -874 135 567
<< psubdiff >>
rect 447 488 507 522
rect 1393 488 1453 522
rect 447 462 481 488
rect 1419 462 1453 488
rect 447 -795 481 -773
rect 1419 -795 1453 -773
rect 447 -829 507 -795
rect 1393 -829 1453 -795
<< nsubdiff >>
rect -907 497 -847 531
rect 39 497 99 531
rect -907 471 -873 497
rect 65 471 99 497
rect -907 -804 -873 -713
rect 65 -804 99 -713
rect -907 -838 -847 -804
rect 39 -838 99 -804
<< psubdiffcont >>
rect 507 488 1393 522
rect 447 -773 481 462
rect 1419 -773 1453 462
rect 507 -829 1393 -795
<< nsubdiffcont >>
rect -847 497 39 531
rect -907 -713 -873 471
rect 65 -713 99 471
rect -847 -838 39 -804
<< poly >>
rect -731 -156 -656 -88
rect -553 -144 -255 -98
rect -151 -154 -79 -88
rect 623 -154 697 -88
rect 865 -144 1035 -98
rect 1277 -150 1307 -86
<< locali >>
rect -907 497 -847 531
rect 39 497 99 531
rect -907 471 -873 497
rect -907 -804 -873 -713
rect 65 471 99 497
rect 65 -804 99 -713
rect -907 -838 -847 -804
rect 39 -838 99 -804
rect 447 488 507 522
rect 1393 488 1453 522
rect 447 462 481 488
rect 447 -795 481 -773
rect 1419 462 1453 488
rect 1419 -795 1453 -773
rect 447 -829 507 -795
rect 1393 -829 1453 -795
<< viali >>
rect -421 497 -387 531
rect -907 -138 -873 -104
rect 65 -138 99 -104
rect -273 -978 -239 -944
<< metal1 >>
rect -433 531 -375 537
rect -433 497 -421 531
rect -387 497 -375 531
rect -433 491 -375 497
rect -421 431 -387 491
rect -388 -37 -387 -7
rect -919 -104 -861 -98
rect -807 -104 -773 -45
rect -719 -94 -685 -41
rect -919 -138 -907 -104
rect -873 -138 -773 -104
rect -919 -144 -861 -138
rect -807 -197 -773 -138
rect -738 -146 -728 -94
rect -676 -146 -666 -94
rect -719 -197 -685 -146
rect -421 -197 -387 -41
rect -123 -95 -89 -41
rect -143 -147 -132 -95
rect -80 -147 -70 -95
rect -35 -104 -1 -45
rect 629 -96 675 -54
rect 53 -104 111 -98
rect -35 -138 65 -104
rect 99 -138 111 -104
rect -123 -197 -89 -147
rect -35 -197 -1 -138
rect 53 -144 111 -138
rect 616 -148 626 -96
rect 678 -148 688 -96
rect 629 -188 675 -148
rect 927 -188 973 -54
rect 1225 -88 1271 -54
rect 1222 -96 1274 -88
rect 1222 -154 1274 -148
rect 1225 -188 1271 -154
rect -273 -938 -239 -732
rect -285 -944 -227 -938
rect -285 -978 -273 -944
rect -239 -978 -227 -944
rect -285 -984 -227 -978
<< via1 >>
rect -728 -146 -676 -94
rect -132 -147 -80 -95
rect 626 -148 678 -96
rect 1222 -148 1274 -96
<< metal2 >>
rect -728 -94 -80 -84
rect -676 -95 -80 -94
rect -676 -146 -132 -95
rect -728 -147 -132 -146
rect 626 -96 678 -86
rect -728 -156 -80 -147
rect 616 -148 626 -96
rect 678 -148 1222 -96
rect 1274 -148 1287 -96
rect 626 -158 678 -148
use sky130_fd_pr__nfet_01v8_8STJTB  sky130_fd_pr__nfet_01v8_8STJTB_1
timestamp 1730520524
transform 1 0 801 0 1 153
box -178 -307 178 307
use sky130_fd_pr__nfet_01v8_8STJTB  sky130_fd_pr__nfet_01v8_8STJTB_2
timestamp 1730520524
transform 1 0 1099 0 1 153
box -178 -307 178 307
use sky130_fd_pr__nfet_01v8_ALPWAK  sky130_fd_pr__nfet_01v8_ALPWAK_1
timestamp 1730520524
transform 1 0 801 0 1 -395
box -178 -307 178 307
use sky130_fd_pr__nfet_01v8_AS47HM  sky130_fd_pr__nfet_01v8_AS47HM_0
timestamp 1730525663
transform 1 0 1099 0 1 -426
box -178 -338 178 338
use sky130_fd_pr__nfet_01v8_LLMDSU  sky130_fd_pr__nfet_01v8_LLMDSU_2
timestamp 1730526150
transform 1 0 608 0 1 153
box -73 -307 73 307
use sky130_fd_pr__nfet_01v8_Q35DSU  sky130_fd_pr__nfet_01v8_Q35DSU_0
timestamp 1730527170
transform 1 0 1292 0 1 184
box -73 -276 73 276
use sky130_fd_pr__nfet_01v8_Q35DSU  sky130_fd_pr__nfet_01v8_Q35DSU_1
timestamp 1730527170
transform 1 0 1292 0 1 -426
box -73 -276 73 276
use sky130_fd_pr__nfet_01v8_Q96DSU  sky130_fd_pr__nfet_01v8_Q96DSU_0
timestamp 1730526150
transform 1 0 608 0 1 -395
box -73 -307 73 307
use sky130_fd_pr__pfet_01v8_D5QVFZ  sky130_fd_pr__pfet_01v8_D5QVFZ_0
timestamp 1730518657
transform 1 0 -255 0 1 157
box -214 -314 214 348
use sky130_fd_pr__pfet_01v8_D5QVFZ  sky130_fd_pr__pfet_01v8_D5QVFZ_1
timestamp 1730518657
transform 1 0 -553 0 1 157
box -214 -314 214 348
use sky130_fd_pr__pfet_01v8_KYWVF3  sky130_fd_pr__pfet_01v8_KYWVF3_0
timestamp 1730525416
transform 1 0 -255 0 1 -435
box -214 -350 214 350
use sky130_fd_pr__pfet_01v8_LL4HGW  sky130_fd_pr__pfet_01v8_LL4HGW_0
timestamp 1730521008
transform 1 0 -746 0 1 -399
box -109 -348 109 314
use sky130_fd_pr__pfet_01v8_LL4HGW  sky130_fd_pr__pfet_01v8_LL4HGW_1
timestamp 1730521008
transform 1 0 -62 0 1 -399
box -109 -348 109 314
use sky130_fd_pr__pfet_01v8_LL49CW  sky130_fd_pr__pfet_01v8_LL49CW_0
timestamp 1730521008
transform 1 0 -746 0 1 157
box -109 -314 109 348
use sky130_fd_pr__pfet_01v8_LL49CW  sky130_fd_pr__pfet_01v8_LL49CW_1
timestamp 1730521008
transform 1 0 -62 0 1 157
box -109 -314 109 348
use sky130_fd_pr__pfet_01v8_UWWVT4  sky130_fd_pr__pfet_01v8_UWWVT4_1
timestamp 1730474680
transform 1 0 -553 0 1 -399
box -214 -348 214 314
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 0 -1 1188 1 0 -1437
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 0 -1 -8 1 0 -1148
box -38 -48 314 592
<< end >>
