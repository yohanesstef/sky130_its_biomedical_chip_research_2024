module freq_psc (clk,
    out,
    rst,
    psc);
 input clk;
 output out;
 input rst;
 input [31:0] psc;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire \counter[0] ;
 wire \counter[10] ;
 wire \counter[11] ;
 wire \counter[12] ;
 wire \counter[13] ;
 wire \counter[14] ;
 wire \counter[15] ;
 wire \counter[16] ;
 wire \counter[17] ;
 wire \counter[18] ;
 wire \counter[19] ;
 wire \counter[1] ;
 wire \counter[20] ;
 wire \counter[21] ;
 wire \counter[22] ;
 wire \counter[23] ;
 wire \counter[24] ;
 wire \counter[25] ;
 wire \counter[26] ;
 wire \counter[27] ;
 wire \counter[28] ;
 wire \counter[29] ;
 wire \counter[2] ;
 wire \counter[30] ;
 wire \counter[31] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \counter[5] ;
 wire \counter[6] ;
 wire \counter[7] ;
 wire \counter[8] ;
 wire \counter[9] ;

 sky130_fd_sc_hd__inv_2 _386_ (.A(\counter[0] ),
    .Y(_066_));
 sky130_fd_sc_hd__inv_2 _387_ (.A(\counter[1] ),
    .Y(_067_));
 sky130_fd_sc_hd__inv_2 _388_ (.A(psc[2]),
    .Y(_068_));
 sky130_fd_sc_hd__inv_2 _389_ (.A(psc[5]),
    .Y(_069_));
 sky130_fd_sc_hd__inv_2 _390_ (.A(psc[6]),
    .Y(_070_));
 sky130_fd_sc_hd__inv_2 _391_ (.A(psc[7]),
    .Y(_071_));
 sky130_fd_sc_hd__inv_2 _392_ (.A(psc[9]),
    .Y(_072_));
 sky130_fd_sc_hd__inv_2 _393_ (.A(\counter[14] ),
    .Y(_073_));
 sky130_fd_sc_hd__inv_2 _394_ (.A(\counter[13] ),
    .Y(_074_));
 sky130_fd_sc_hd__inv_2 _395_ (.A(\counter[12] ),
    .Y(_075_));
 sky130_fd_sc_hd__inv_2 _396_ (.A(\counter[10] ),
    .Y(_076_));
 sky130_fd_sc_hd__inv_2 _397_ (.A(\counter[9] ),
    .Y(_077_));
 sky130_fd_sc_hd__inv_2 _398_ (.A(psc[29]),
    .Y(_078_));
 sky130_fd_sc_hd__inv_2 _399_ (.A(psc[28]),
    .Y(_079_));
 sky130_fd_sc_hd__inv_2 _400_ (.A(psc[26]),
    .Y(_080_));
 sky130_fd_sc_hd__inv_2 _401_ (.A(psc[25]),
    .Y(_081_));
 sky130_fd_sc_hd__inv_2 _402_ (.A(psc[24]),
    .Y(_082_));
 sky130_fd_sc_hd__inv_2 _403_ (.A(psc[23]),
    .Y(_083_));
 sky130_fd_sc_hd__inv_2 _404_ (.A(psc[22]),
    .Y(_084_));
 sky130_fd_sc_hd__inv_2 _405_ (.A(psc[21]),
    .Y(_085_));
 sky130_fd_sc_hd__inv_2 _406_ (.A(psc[19]),
    .Y(_086_));
 sky130_fd_sc_hd__inv_2 _407_ (.A(psc[18]),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _408_ (.A(psc[17]),
    .Y(_088_));
 sky130_fd_sc_hd__inv_2 _409_ (.A(psc[16]),
    .Y(_089_));
 sky130_fd_sc_hd__inv_2 _410_ (.A(psc[30]),
    .Y(_090_));
 sky130_fd_sc_hd__inv_2 _411_ (.A(psc[31]),
    .Y(_091_));
 sky130_fd_sc_hd__inv_2 _412_ (.A(\counter[30] ),
    .Y(_092_));
 sky130_fd_sc_hd__inv_2 _413_ (.A(\counter[27] ),
    .Y(_093_));
 sky130_fd_sc_hd__inv_2 _414_ (.A(\counter[26] ),
    .Y(_094_));
 sky130_fd_sc_hd__inv_2 _415_ (.A(rst),
    .Y(_033_));
 sky130_fd_sc_hd__or2_2 _416_ (.A(psc[0]),
    .B(psc[1]),
    .X(_095_));
 sky130_fd_sc_hd__or3_2 _417_ (.A(psc[0]),
    .B(psc[1]),
    .C(psc[2]),
    .X(_096_));
 sky130_fd_sc_hd__or4_2 _418_ (.A(psc[0]),
    .B(psc[1]),
    .C(psc[2]),
    .D(psc[3]),
    .X(_097_));
 sky130_fd_sc_hd__nor2_2 _419_ (.A(psc[4]),
    .B(_097_),
    .Y(_098_));
 sky130_fd_sc_hd__or4_2 _420_ (.A(psc[5]),
    .B(psc[4]),
    .C(psc[6]),
    .D(_097_),
    .X(_099_));
 sky130_fd_sc_hd__or3_2 _421_ (.A(psc[7]),
    .B(psc[8]),
    .C(_099_),
    .X(_100_));
 sky130_fd_sc_hd__or4_2 _422_ (.A(psc[7]),
    .B(psc[9]),
    .C(psc[8]),
    .D(_099_),
    .X(_101_));
 sky130_fd_sc_hd__or3_2 _423_ (.A(psc[10]),
    .B(psc[9]),
    .C(psc[8]),
    .X(_102_));
 sky130_fd_sc_hd__or4_2 _424_ (.A(psc[7]),
    .B(psc[11]),
    .C(_099_),
    .D(_102_),
    .X(_103_));
 sky130_fd_sc_hd__or2_2 _425_ (.A(psc[13]),
    .B(psc[12]),
    .X(_104_));
 sky130_fd_sc_hd__nor2_2 _426_ (.A(_103_),
    .B(_104_),
    .Y(_105_));
 sky130_fd_sc_hd__nor4_2 _427_ (.A(psc[14]),
    .B(psc[15]),
    .C(_103_),
    .D(_104_),
    .Y(_106_));
 sky130_fd_sc_hd__or4_2 _428_ (.A(psc[14]),
    .B(psc[15]),
    .C(_103_),
    .D(_104_),
    .X(_107_));
 sky130_fd_sc_hd__or4_2 _429_ (.A(psc[23]),
    .B(psc[20]),
    .C(psc[19]),
    .D(psc[16]),
    .X(_108_));
 sky130_fd_sc_hd__or2_2 _430_ (.A(psc[18]),
    .B(psc[17]),
    .X(_109_));
 sky130_fd_sc_hd__or4_2 _431_ (.A(psc[22]),
    .B(psc[21]),
    .C(_108_),
    .D(_109_),
    .X(_110_));
 sky130_fd_sc_hd__inv_2 _432_ (.A(_110_),
    .Y(_111_));
 sky130_fd_sc_hd__nor2_2 _433_ (.A(psc[20]),
    .B(psc[19]),
    .Y(_112_));
 sky130_fd_sc_hd__nand2_2 _434_ (.A(_106_),
    .B(_111_),
    .Y(_113_));
 sky130_fd_sc_hd__or4_2 _435_ (.A(psc[25]),
    .B(psc[24]),
    .C(_107_),
    .D(_110_),
    .X(_114_));
 sky130_fd_sc_hd__and4b_2 _436_ (.A_N(psc[27]),
    .B(_080_),
    .C(_081_),
    .D(_082_),
    .X(_115_));
 sky130_fd_sc_hd__or3_2 _437_ (.A(psc[27]),
    .B(psc[26]),
    .C(_114_),
    .X(_116_));
 sky130_fd_sc_hd__or4b_2 _438_ (.A(psc[28]),
    .B(_107_),
    .C(_110_),
    .D_N(_115_),
    .X(_117_));
 sky130_fd_sc_hd__or3_2 _439_ (.A(psc[29]),
    .B(psc[30]),
    .C(_117_),
    .X(_118_));
 sky130_fd_sc_hd__o31ai_2 _440_ (.A1(psc[29]),
    .A2(psc[30]),
    .A3(_117_),
    .B1(psc[31]),
    .Y(_119_));
 sky130_fd_sc_hd__or4_2 _441_ (.A(psc[29]),
    .B(psc[30]),
    .C(psc[31]),
    .D(_117_),
    .X(_120_));
 sky130_fd_sc_hd__a21oi_2 _442_ (.A1(_119_),
    .A2(_120_),
    .B1(\counter[31] ),
    .Y(_121_));
 sky130_fd_sc_hd__o21ai_2 _443_ (.A1(psc[29]),
    .A2(_117_),
    .B1(psc[30]),
    .Y(_122_));
 sky130_fd_sc_hd__and3_2 _444_ (.A(\counter[30] ),
    .B(_118_),
    .C(_122_),
    .X(_123_));
 sky130_fd_sc_hd__a31oi_2 _445_ (.A1(\counter[31] ),
    .A2(_119_),
    .A3(_120_),
    .B1(_123_),
    .Y(_124_));
 sky130_fd_sc_hd__xnor2_2 _446_ (.A(_078_),
    .B(_117_),
    .Y(_125_));
 sky130_fd_sc_hd__a31o_2 _447_ (.A1(_106_),
    .A2(_111_),
    .A3(_115_),
    .B1(_079_),
    .X(_126_));
 sky130_fd_sc_hd__and3_2 _448_ (.A(\counter[28] ),
    .B(_117_),
    .C(_126_),
    .X(_127_));
 sky130_fd_sc_hd__a21oi_2 _449_ (.A1(\counter[29] ),
    .A2(_125_),
    .B1(_127_),
    .Y(_128_));
 sky130_fd_sc_hd__nor2_2 _450_ (.A(\counter[29] ),
    .B(_125_),
    .Y(_129_));
 sky130_fd_sc_hd__a21oi_2 _451_ (.A1(_118_),
    .A2(_122_),
    .B1(\counter[30] ),
    .Y(_130_));
 sky130_fd_sc_hd__o31a_2 _452_ (.A1(_128_),
    .A2(_129_),
    .A3(_130_),
    .B1(_124_),
    .X(_131_));
 sky130_fd_sc_hd__a21oi_2 _453_ (.A1(_117_),
    .A2(_126_),
    .B1(\counter[28] ),
    .Y(_132_));
 sky130_fd_sc_hd__a211o_2 _454_ (.A1(\counter[29] ),
    .A2(_125_),
    .B1(_127_),
    .C1(_132_),
    .X(_133_));
 sky130_fd_sc_hd__nor4_2 _455_ (.A(_121_),
    .B(_129_),
    .C(_130_),
    .D(_133_),
    .Y(_134_));
 sky130_fd_sc_hd__and2_2 _456_ (.A(_124_),
    .B(_134_),
    .X(_135_));
 sky130_fd_sc_hd__a31o_2 _457_ (.A1(_082_),
    .A2(_106_),
    .A3(_111_),
    .B1(_081_),
    .X(_136_));
 sky130_fd_sc_hd__and2_2 _458_ (.A(_114_),
    .B(_136_),
    .X(_137_));
 sky130_fd_sc_hd__xnor2_2 _459_ (.A(_082_),
    .B(_113_),
    .Y(_138_));
 sky130_fd_sc_hd__a22o_2 _460_ (.A1(\counter[25] ),
    .A2(_137_),
    .B1(_138_),
    .B2(\counter[24] ),
    .X(_139_));
 sky130_fd_sc_hd__o21ai_2 _461_ (.A1(psc[26]),
    .A2(_114_),
    .B1(psc[27]),
    .Y(_140_));
 sky130_fd_sc_hd__a21o_2 _462_ (.A1(_116_),
    .A2(_140_),
    .B1(\counter[27] ),
    .X(_141_));
 sky130_fd_sc_hd__xnor2_2 _463_ (.A(_080_),
    .B(_114_),
    .Y(_142_));
 sky130_fd_sc_hd__nand2_2 _464_ (.A(\counter[26] ),
    .B(_142_),
    .Y(_143_));
 sky130_fd_sc_hd__or2_2 _465_ (.A(\counter[26] ),
    .B(_142_),
    .X(_144_));
 sky130_fd_sc_hd__or2_2 _466_ (.A(\counter[25] ),
    .B(_137_),
    .X(_145_));
 sky130_fd_sc_hd__and4_2 _467_ (.A(_141_),
    .B(_143_),
    .C(_144_),
    .D(_145_),
    .X(_146_));
 sky130_fd_sc_hd__and3_2 _468_ (.A(_141_),
    .B(_143_),
    .C(_144_),
    .X(_147_));
 sky130_fd_sc_hd__and3_2 _469_ (.A(\counter[27] ),
    .B(_116_),
    .C(_140_),
    .X(_148_));
 sky130_fd_sc_hd__and3_2 _470_ (.A(\counter[26] ),
    .B(_141_),
    .C(_142_),
    .X(_149_));
 sky130_fd_sc_hd__a211o_2 _471_ (.A1(_139_),
    .A2(_146_),
    .B1(_148_),
    .C1(_149_),
    .X(_150_));
 sky130_fd_sc_hd__o2bb2a_2 _472_ (.A1_N(_135_),
    .A2_N(_150_),
    .B1(_121_),
    .B2(_131_),
    .X(_151_));
 sky130_fd_sc_hd__and3b_2 _473_ (.A_N(_109_),
    .B(_089_),
    .C(_106_),
    .X(_152_));
 sky130_fd_sc_hd__and4b_2 _474_ (.A_N(_109_),
    .B(_089_),
    .C(_106_),
    .D(_112_),
    .X(_153_));
 sky130_fd_sc_hd__or3b_2 _475_ (.A(psc[22]),
    .B(psc[21]),
    .C_N(_153_),
    .X(_154_));
 sky130_fd_sc_hd__a31o_2 _476_ (.A1(_084_),
    .A2(_085_),
    .A3(_153_),
    .B1(_083_),
    .X(_155_));
 sky130_fd_sc_hd__and3_2 _477_ (.A(\counter[23] ),
    .B(_113_),
    .C(_155_),
    .X(_156_));
 sky130_fd_sc_hd__a21o_2 _478_ (.A1(_085_),
    .A2(_153_),
    .B1(_084_),
    .X(_157_));
 sky130_fd_sc_hd__a31o_2 _479_ (.A1(\counter[22] ),
    .A2(_154_),
    .A3(_157_),
    .B1(_156_),
    .X(_158_));
 sky130_fd_sc_hd__a21o_2 _480_ (.A1(_113_),
    .A2(_155_),
    .B1(\counter[23] ),
    .X(_159_));
 sky130_fd_sc_hd__xnor2_2 _481_ (.A(psc[21]),
    .B(_153_),
    .Y(_160_));
 sky130_fd_sc_hd__a21o_2 _482_ (.A1(_154_),
    .A2(_157_),
    .B1(\counter[22] ),
    .X(_161_));
 sky130_fd_sc_hd__o211ai_2 _483_ (.A1(\counter[21] ),
    .A2(_160_),
    .B1(_161_),
    .C1(_159_),
    .Y(_162_));
 sky130_fd_sc_hd__o41a_2 _484_ (.A1(psc[19]),
    .A2(psc[16]),
    .A3(_107_),
    .A4(_109_),
    .B1(psc[20]),
    .X(_163_));
 sky130_fd_sc_hd__nor2_2 _485_ (.A(_153_),
    .B(_163_),
    .Y(_164_));
 sky130_fd_sc_hd__a22oi_2 _486_ (.A1(\counter[21] ),
    .A2(_160_),
    .B1(_164_),
    .B2(\counter[20] ),
    .Y(_165_));
 sky130_fd_sc_hd__o21ai_2 _487_ (.A1(\counter[20] ),
    .A2(_164_),
    .B1(_165_),
    .Y(_166_));
 sky130_fd_sc_hd__xnor2_2 _488_ (.A(psc[19]),
    .B(_152_),
    .Y(_167_));
 sky130_fd_sc_hd__or3_2 _489_ (.A(psc[17]),
    .B(psc[16]),
    .C(_107_),
    .X(_168_));
 sky130_fd_sc_hd__a21oi_2 _490_ (.A1(psc[18]),
    .A2(_168_),
    .B1(_152_),
    .Y(_169_));
 sky130_fd_sc_hd__a22o_2 _491_ (.A1(\counter[19] ),
    .A2(_167_),
    .B1(_169_),
    .B2(\counter[18] ),
    .X(_170_));
 sky130_fd_sc_hd__o21a_2 _492_ (.A1(\counter[19] ),
    .A2(_167_),
    .B1(_170_),
    .X(_171_));
 sky130_fd_sc_hd__o22a_2 _493_ (.A1(\counter[19] ),
    .A2(_167_),
    .B1(_169_),
    .B2(\counter[18] ),
    .X(_172_));
 sky130_fd_sc_hd__a21o_2 _494_ (.A1(_089_),
    .A2(_106_),
    .B1(_088_),
    .X(_173_));
 sky130_fd_sc_hd__and2_2 _495_ (.A(_168_),
    .B(_173_),
    .X(_174_));
 sky130_fd_sc_hd__nor2_2 _496_ (.A(\counter[17] ),
    .B(_174_),
    .Y(_175_));
 sky130_fd_sc_hd__xnor2_2 _497_ (.A(psc[16]),
    .B(_106_),
    .Y(_176_));
 sky130_fd_sc_hd__a22o_2 _498_ (.A1(\counter[17] ),
    .A2(_174_),
    .B1(_176_),
    .B2(\counter[16] ),
    .X(_177_));
 sky130_fd_sc_hd__and3b_2 _499_ (.A_N(_175_),
    .B(_177_),
    .C(_172_),
    .X(_178_));
 sky130_fd_sc_hd__nor2_2 _500_ (.A(_171_),
    .B(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__o31a_2 _501_ (.A1(psc[14]),
    .A2(_103_),
    .A3(_104_),
    .B1(psc[15]),
    .X(_180_));
 sky130_fd_sc_hd__nor2_2 _502_ (.A(_106_),
    .B(_180_),
    .Y(_181_));
 sky130_fd_sc_hd__xnor2_2 _503_ (.A(psc[14]),
    .B(_105_),
    .Y(_182_));
 sky130_fd_sc_hd__a22o_2 _504_ (.A1(\counter[15] ),
    .A2(_181_),
    .B1(_182_),
    .B2(\counter[14] ),
    .X(_183_));
 sky130_fd_sc_hd__or2_2 _505_ (.A(psc[12]),
    .B(_103_),
    .X(_184_));
 sky130_fd_sc_hd__a21oi_2 _506_ (.A1(psc[13]),
    .A2(_184_),
    .B1(_105_),
    .Y(_185_));
 sky130_fd_sc_hd__o22a_2 _507_ (.A1(\counter[14] ),
    .A2(_182_),
    .B1(_185_),
    .B2(\counter[13] ),
    .X(_186_));
 sky130_fd_sc_hd__nand2_2 _508_ (.A(psc[12]),
    .B(_103_),
    .Y(_187_));
 sky130_fd_sc_hd__and2_2 _509_ (.A(_184_),
    .B(_187_),
    .X(_188_));
 sky130_fd_sc_hd__a22o_2 _510_ (.A1(\counter[13] ),
    .A2(_185_),
    .B1(_188_),
    .B2(\counter[12] ),
    .X(_189_));
 sky130_fd_sc_hd__o21ai_2 _511_ (.A1(psc[10]),
    .A2(_101_),
    .B1(psc[11]),
    .Y(_190_));
 sky130_fd_sc_hd__and2_2 _512_ (.A(_103_),
    .B(_190_),
    .X(_191_));
 sky130_fd_sc_hd__xor2_2 _513_ (.A(psc[10]),
    .B(_101_),
    .X(_192_));
 sky130_fd_sc_hd__xnor2_2 _514_ (.A(_072_),
    .B(_100_),
    .Y(_193_));
 sky130_fd_sc_hd__a22o_2 _515_ (.A1(\counter[10] ),
    .A2(_192_),
    .B1(_193_),
    .B2(\counter[9] ),
    .X(_194_));
 sky130_fd_sc_hd__or2_2 _516_ (.A(\counter[9] ),
    .B(_193_),
    .X(_195_));
 sky130_fd_sc_hd__o21ai_2 _517_ (.A1(psc[7]),
    .A2(_099_),
    .B1(psc[8]),
    .Y(_196_));
 sky130_fd_sc_hd__and2_2 _518_ (.A(_100_),
    .B(_196_),
    .X(_197_));
 sky130_fd_sc_hd__xnor2_2 _519_ (.A(_071_),
    .B(_099_),
    .Y(_198_));
 sky130_fd_sc_hd__nand2_2 _520_ (.A(psc[3]),
    .B(_096_),
    .Y(_199_));
 sky130_fd_sc_hd__and2_2 _521_ (.A(_097_),
    .B(_199_),
    .X(_200_));
 sky130_fd_sc_hd__nand2_2 _522_ (.A(psc[2]),
    .B(_095_),
    .Y(_201_));
 sky130_fd_sc_hd__a21o_2 _523_ (.A1(_096_),
    .A2(_201_),
    .B1(\counter[2] ),
    .X(_202_));
 sky130_fd_sc_hd__and3_2 _524_ (.A(\counter[2] ),
    .B(_096_),
    .C(_201_),
    .X(_203_));
 sky130_fd_sc_hd__nand2_2 _525_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .Y(_204_));
 sky130_fd_sc_hd__o211ai_2 _526_ (.A1(psc[0]),
    .A2(_066_),
    .B1(psc[1]),
    .C1(_067_),
    .Y(_205_));
 sky130_fd_sc_hd__a21bo_2 _527_ (.A1(_095_),
    .A2(_205_),
    .B1_N(_204_),
    .X(_206_));
 sky130_fd_sc_hd__a221o_2 _528_ (.A1(\counter[3] ),
    .A2(_200_),
    .B1(_202_),
    .B2(_206_),
    .C1(_203_),
    .X(_207_));
 sky130_fd_sc_hd__nand2_2 _529_ (.A(psc[4]),
    .B(_097_),
    .Y(_208_));
 sky130_fd_sc_hd__and2b_2 _530_ (.A_N(_098_),
    .B(_208_),
    .X(_209_));
 sky130_fd_sc_hd__o221a_2 _531_ (.A1(\counter[3] ),
    .A2(_200_),
    .B1(_209_),
    .B2(\counter[4] ),
    .C1(_207_),
    .X(_210_));
 sky130_fd_sc_hd__xnor2_2 _532_ (.A(psc[5]),
    .B(_098_),
    .Y(_211_));
 sky130_fd_sc_hd__a22o_2 _533_ (.A1(\counter[4] ),
    .A2(_209_),
    .B1(_211_),
    .B2(\counter[5] ),
    .X(_212_));
 sky130_fd_sc_hd__a21o_2 _534_ (.A1(_069_),
    .A2(_098_),
    .B1(_070_),
    .X(_213_));
 sky130_fd_sc_hd__and2_2 _535_ (.A(_099_),
    .B(_213_),
    .X(_214_));
 sky130_fd_sc_hd__or2_2 _536_ (.A(\counter[6] ),
    .B(_214_),
    .X(_215_));
 sky130_fd_sc_hd__o221a_2 _537_ (.A1(\counter[5] ),
    .A2(_211_),
    .B1(_212_),
    .B2(_210_),
    .C1(_215_),
    .X(_216_));
 sky130_fd_sc_hd__a22o_2 _538_ (.A1(\counter[7] ),
    .A2(_198_),
    .B1(_214_),
    .B2(\counter[6] ),
    .X(_217_));
 sky130_fd_sc_hd__o22a_2 _539_ (.A1(\counter[11] ),
    .A2(_191_),
    .B1(_192_),
    .B2(\counter[10] ),
    .X(_218_));
 sky130_fd_sc_hd__a31o_2 _540_ (.A1(\counter[8] ),
    .A2(_195_),
    .A3(_197_),
    .B1(_194_),
    .X(_219_));
 sky130_fd_sc_hd__a22o_2 _541_ (.A1(\counter[11] ),
    .A2(_191_),
    .B1(_218_),
    .B2(_219_),
    .X(_220_));
 sky130_fd_sc_hd__o2bb2a_2 _542_ (.A1_N(\counter[8] ),
    .A2_N(_197_),
    .B1(_193_),
    .B2(\counter[9] ),
    .X(_221_));
 sky130_fd_sc_hd__o221a_2 _543_ (.A1(\counter[8] ),
    .A2(_197_),
    .B1(_198_),
    .B2(\counter[7] ),
    .C1(_221_),
    .X(_222_));
 sky130_fd_sc_hd__o21ba_2 _544_ (.A1(_216_),
    .A2(_217_),
    .B1_N(_194_),
    .X(_223_));
 sky130_fd_sc_hd__a31o_2 _545_ (.A1(_218_),
    .A2(_222_),
    .A3(_223_),
    .B1(_220_),
    .X(_224_));
 sky130_fd_sc_hd__nor2_2 _546_ (.A(\counter[16] ),
    .B(_176_),
    .Y(_225_));
 sky130_fd_sc_hd__or3_2 _547_ (.A(_158_),
    .B(_162_),
    .C(_166_),
    .X(_226_));
 sky130_fd_sc_hd__or3_2 _548_ (.A(_158_),
    .B(_162_),
    .C(_165_),
    .X(_227_));
 sky130_fd_sc_hd__nand2_2 _549_ (.A(_158_),
    .B(_159_),
    .Y(_228_));
 sky130_fd_sc_hd__or2_2 _550_ (.A(\counter[24] ),
    .B(_138_),
    .X(_229_));
 sky130_fd_sc_hd__and3b_2 _551_ (.A_N(_139_),
    .B(_145_),
    .C(_229_),
    .X(_230_));
 sky130_fd_sc_hd__nand4_2 _552_ (.A(_124_),
    .B(_134_),
    .C(_147_),
    .D(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__or2_2 _553_ (.A(_148_),
    .B(_231_),
    .X(_232_));
 sky130_fd_sc_hd__nor2_2 _554_ (.A(_183_),
    .B(_189_),
    .Y(_233_));
 sky130_fd_sc_hd__o221a_2 _555_ (.A1(\counter[15] ),
    .A2(_181_),
    .B1(_188_),
    .B2(\counter[12] ),
    .C1(_186_),
    .X(_234_));
 sky130_fd_sc_hd__a21o_2 _556_ (.A1(_186_),
    .A2(_189_),
    .B1(_183_),
    .X(_235_));
 sky130_fd_sc_hd__o21a_2 _557_ (.A1(\counter[15] ),
    .A2(_181_),
    .B1(_235_),
    .X(_236_));
 sky130_fd_sc_hd__a31oi_2 _558_ (.A1(_224_),
    .A2(_233_),
    .A3(_234_),
    .B1(_236_),
    .Y(_237_));
 sky130_fd_sc_hd__a221o_2 _559_ (.A1(\counter[19] ),
    .A2(_167_),
    .B1(_169_),
    .B2(\counter[18] ),
    .C1(_225_),
    .X(_238_));
 sky130_fd_sc_hd__or4b_2 _560_ (.A(_175_),
    .B(_177_),
    .C(_238_),
    .D_N(_172_),
    .X(_239_));
 sky130_fd_sc_hd__or4_2 _561_ (.A(_158_),
    .B(_162_),
    .C(_166_),
    .D(_239_),
    .X(_240_));
 sky130_fd_sc_hd__or4_2 _562_ (.A(_148_),
    .B(_231_),
    .C(_237_),
    .D(_240_),
    .X(_241_));
 sky130_fd_sc_hd__o211a_2 _563_ (.A1(_179_),
    .A2(_226_),
    .B1(_227_),
    .C1(_228_),
    .X(_242_));
 sky130_fd_sc_hd__o211a_2 _564_ (.A1(_232_),
    .A2(_242_),
    .B1(_241_),
    .C1(_151_),
    .X(_243_));
 sky130_fd_sc_hd__and2_2 _565_ (.A(_066_),
    .B(_243_),
    .X(_000_));
 sky130_fd_sc_hd__or2_2 _566_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .X(_244_));
 sky130_fd_sc_hd__and3_2 _567_ (.A(_204_),
    .B(_243_),
    .C(_244_),
    .X(_011_));
 sky130_fd_sc_hd__and3_2 _568_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .C(\counter[2] ),
    .X(_245_));
 sky130_fd_sc_hd__a21o_2 _569_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .B1(\counter[2] ),
    .X(_246_));
 sky130_fd_sc_hd__and3b_2 _570_ (.A_N(_245_),
    .B(_246_),
    .C(_243_),
    .X(_022_));
 sky130_fd_sc_hd__and4_2 _571_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .C(\counter[3] ),
    .D(\counter[2] ),
    .X(_247_));
 sky130_fd_sc_hd__or2_2 _572_ (.A(\counter[3] ),
    .B(_245_),
    .X(_248_));
 sky130_fd_sc_hd__and3b_2 _573_ (.A_N(_247_),
    .B(_248_),
    .C(_243_),
    .X(_025_));
 sky130_fd_sc_hd__nand2_2 _574_ (.A(\counter[4] ),
    .B(_247_),
    .Y(_249_));
 sky130_fd_sc_hd__or2_2 _575_ (.A(\counter[4] ),
    .B(_247_),
    .X(_250_));
 sky130_fd_sc_hd__and3_2 _576_ (.A(_243_),
    .B(_249_),
    .C(_250_),
    .X(_026_));
 sky130_fd_sc_hd__and3_2 _577_ (.A(\counter[5] ),
    .B(\counter[4] ),
    .C(_247_),
    .X(_251_));
 sky130_fd_sc_hd__a21o_2 _578_ (.A1(\counter[4] ),
    .A2(_247_),
    .B1(\counter[5] ),
    .X(_252_));
 sky130_fd_sc_hd__and3b_2 _579_ (.A_N(_251_),
    .B(_252_),
    .C(_243_),
    .X(_027_));
 sky130_fd_sc_hd__and4_2 _580_ (.A(\counter[6] ),
    .B(\counter[5] ),
    .C(\counter[4] ),
    .D(_247_),
    .X(_253_));
 sky130_fd_sc_hd__or2_2 _581_ (.A(\counter[6] ),
    .B(_251_),
    .X(_254_));
 sky130_fd_sc_hd__and3b_2 _582_ (.A_N(_253_),
    .B(_254_),
    .C(_243_),
    .X(_028_));
 sky130_fd_sc_hd__and2_2 _583_ (.A(\counter[7] ),
    .B(_253_),
    .X(_255_));
 sky130_fd_sc_hd__or2_2 _584_ (.A(\counter[7] ),
    .B(_253_),
    .X(_256_));
 sky130_fd_sc_hd__and3b_2 _585_ (.A_N(_255_),
    .B(_256_),
    .C(_243_),
    .X(_029_));
 sky130_fd_sc_hd__nand2_2 _586_ (.A(\counter[8] ),
    .B(_255_),
    .Y(_257_));
 sky130_fd_sc_hd__or2_2 _587_ (.A(\counter[8] ),
    .B(_255_),
    .X(_258_));
 sky130_fd_sc_hd__and3_2 _588_ (.A(_243_),
    .B(_257_),
    .C(_258_),
    .X(_030_));
 sky130_fd_sc_hd__nand2_2 _589_ (.A(_077_),
    .B(_257_),
    .Y(_259_));
 sky130_fd_sc_hd__and2_2 _590_ (.A(\counter[9] ),
    .B(\counter[8] ),
    .X(_260_));
 sky130_fd_sc_hd__and3_2 _591_ (.A(\counter[7] ),
    .B(_253_),
    .C(_260_),
    .X(_261_));
 sky130_fd_sc_hd__and3b_2 _592_ (.A_N(_261_),
    .B(_243_),
    .C(_259_),
    .X(_031_));
 sky130_fd_sc_hd__and4_2 _593_ (.A(\counter[7] ),
    .B(\counter[10] ),
    .C(_253_),
    .D(_260_),
    .X(_262_));
 sky130_fd_sc_hd__or2_2 _594_ (.A(\counter[10] ),
    .B(_261_),
    .X(_263_));
 sky130_fd_sc_hd__and3b_2 _595_ (.A_N(_262_),
    .B(_263_),
    .C(_243_),
    .X(_001_));
 sky130_fd_sc_hd__or2_2 _596_ (.A(\counter[11] ),
    .B(_262_),
    .X(_264_));
 sky130_fd_sc_hd__and2_2 _597_ (.A(\counter[11] ),
    .B(_262_),
    .X(_265_));
 sky130_fd_sc_hd__and3b_2 _598_ (.A_N(_265_),
    .B(_243_),
    .C(_264_),
    .X(_002_));
 sky130_fd_sc_hd__or2_2 _599_ (.A(\counter[12] ),
    .B(_265_),
    .X(_266_));
 sky130_fd_sc_hd__and3_2 _600_ (.A(\counter[12] ),
    .B(\counter[11] ),
    .C(_262_),
    .X(_267_));
 sky130_fd_sc_hd__and3b_2 _601_ (.A_N(_267_),
    .B(_243_),
    .C(_266_),
    .X(_003_));
 sky130_fd_sc_hd__or2_2 _602_ (.A(\counter[13] ),
    .B(_267_),
    .X(_268_));
 sky130_fd_sc_hd__and4_2 _603_ (.A(\counter[13] ),
    .B(\counter[12] ),
    .C(\counter[11] ),
    .D(_262_),
    .X(_269_));
 sky130_fd_sc_hd__and3b_2 _604_ (.A_N(_269_),
    .B(_243_),
    .C(_268_),
    .X(_004_));
 sky130_fd_sc_hd__nand2_2 _605_ (.A(\counter[14] ),
    .B(_269_),
    .Y(_270_));
 sky130_fd_sc_hd__or2_2 _606_ (.A(\counter[14] ),
    .B(_269_),
    .X(_271_));
 sky130_fd_sc_hd__and3_2 _607_ (.A(_243_),
    .B(_270_),
    .C(_271_),
    .X(_005_));
 sky130_fd_sc_hd__a21o_2 _608_ (.A1(\counter[14] ),
    .A2(_269_),
    .B1(\counter[15] ),
    .X(_272_));
 sky130_fd_sc_hd__and3_2 _609_ (.A(\counter[15] ),
    .B(\counter[14] ),
    .C(_269_),
    .X(_273_));
 sky130_fd_sc_hd__and3b_2 _610_ (.A_N(_273_),
    .B(_243_),
    .C(_272_),
    .X(_006_));
 sky130_fd_sc_hd__and2_2 _611_ (.A(\counter[16] ),
    .B(_273_),
    .X(_274_));
 sky130_fd_sc_hd__or2_2 _612_ (.A(\counter[16] ),
    .B(_273_),
    .X(_275_));
 sky130_fd_sc_hd__and3b_2 _613_ (.A_N(_274_),
    .B(_275_),
    .C(_243_),
    .X(_007_));
 sky130_fd_sc_hd__and2_2 _614_ (.A(\counter[17] ),
    .B(\counter[16] ),
    .X(_276_));
 sky130_fd_sc_hd__and4_2 _615_ (.A(\counter[15] ),
    .B(\counter[14] ),
    .C(_269_),
    .D(_276_),
    .X(_277_));
 sky130_fd_sc_hd__inv_2 _616_ (.A(_277_),
    .Y(_278_));
 sky130_fd_sc_hd__o211a_2 _617_ (.A1(\counter[17] ),
    .A2(_274_),
    .B1(_278_),
    .C1(_243_),
    .X(_008_));
 sky130_fd_sc_hd__and2_2 _618_ (.A(\counter[18] ),
    .B(_277_),
    .X(_279_));
 sky130_fd_sc_hd__or2_2 _619_ (.A(\counter[18] ),
    .B(_277_),
    .X(_280_));
 sky130_fd_sc_hd__and3b_2 _620_ (.A_N(_279_),
    .B(_280_),
    .C(_243_),
    .X(_009_));
 sky130_fd_sc_hd__or2_2 _621_ (.A(\counter[19] ),
    .B(_279_),
    .X(_281_));
 sky130_fd_sc_hd__and3_2 _622_ (.A(\counter[19] ),
    .B(\counter[18] ),
    .C(_277_),
    .X(_282_));
 sky130_fd_sc_hd__and3b_2 _623_ (.A_N(_282_),
    .B(_243_),
    .C(_281_),
    .X(_010_));
 sky130_fd_sc_hd__and4_2 _624_ (.A(\counter[20] ),
    .B(\counter[19] ),
    .C(\counter[18] ),
    .D(_277_),
    .X(_283_));
 sky130_fd_sc_hd__or2_2 _625_ (.A(\counter[20] ),
    .B(_282_),
    .X(_284_));
 sky130_fd_sc_hd__and3b_2 _626_ (.A_N(_283_),
    .B(_284_),
    .C(_243_),
    .X(_012_));
 sky130_fd_sc_hd__or2_2 _627_ (.A(\counter[21] ),
    .B(_283_),
    .X(_285_));
 sky130_fd_sc_hd__nand2_2 _628_ (.A(\counter[21] ),
    .B(_283_),
    .Y(_286_));
 sky130_fd_sc_hd__and3_2 _629_ (.A(_243_),
    .B(_285_),
    .C(_286_),
    .X(_013_));
 sky130_fd_sc_hd__and3_2 _630_ (.A(\counter[22] ),
    .B(\counter[21] ),
    .C(_283_),
    .X(_287_));
 sky130_fd_sc_hd__a21o_2 _631_ (.A1(\counter[21] ),
    .A2(_283_),
    .B1(\counter[22] ),
    .X(_288_));
 sky130_fd_sc_hd__and3b_2 _632_ (.A_N(_287_),
    .B(_288_),
    .C(_243_),
    .X(_014_));
 sky130_fd_sc_hd__or2_2 _633_ (.A(\counter[23] ),
    .B(_287_),
    .X(_289_));
 sky130_fd_sc_hd__and4_2 _634_ (.A(\counter[23] ),
    .B(\counter[22] ),
    .C(\counter[21] ),
    .D(_283_),
    .X(_290_));
 sky130_fd_sc_hd__and3b_2 _635_ (.A_N(_290_),
    .B(_243_),
    .C(_289_),
    .X(_015_));
 sky130_fd_sc_hd__nand2_2 _636_ (.A(\counter[24] ),
    .B(_290_),
    .Y(_291_));
 sky130_fd_sc_hd__or2_2 _637_ (.A(\counter[24] ),
    .B(_290_),
    .X(_292_));
 sky130_fd_sc_hd__and3_2 _638_ (.A(_243_),
    .B(_291_),
    .C(_292_),
    .X(_016_));
 sky130_fd_sc_hd__a21o_2 _639_ (.A1(\counter[24] ),
    .A2(_290_),
    .B1(\counter[25] ),
    .X(_293_));
 sky130_fd_sc_hd__and3_2 _640_ (.A(\counter[25] ),
    .B(\counter[24] ),
    .C(_290_),
    .X(_294_));
 sky130_fd_sc_hd__and3b_2 _641_ (.A_N(_294_),
    .B(_243_),
    .C(_293_),
    .X(_017_));
 sky130_fd_sc_hd__and4_2 _642_ (.A(\counter[26] ),
    .B(\counter[25] ),
    .C(\counter[24] ),
    .D(_290_),
    .X(_295_));
 sky130_fd_sc_hd__or2_2 _643_ (.A(\counter[26] ),
    .B(_294_),
    .X(_296_));
 sky130_fd_sc_hd__and3b_2 _644_ (.A_N(_295_),
    .B(_296_),
    .C(_243_),
    .X(_018_));
 sky130_fd_sc_hd__or2_2 _645_ (.A(\counter[27] ),
    .B(_295_),
    .X(_297_));
 sky130_fd_sc_hd__nand2_2 _646_ (.A(\counter[27] ),
    .B(_295_),
    .Y(_298_));
 sky130_fd_sc_hd__and3_2 _647_ (.A(_243_),
    .B(_297_),
    .C(_298_),
    .X(_019_));
 sky130_fd_sc_hd__and3_2 _648_ (.A(\counter[28] ),
    .B(\counter[27] ),
    .C(_295_),
    .X(_299_));
 sky130_fd_sc_hd__a21o_2 _649_ (.A1(\counter[27] ),
    .A2(_295_),
    .B1(\counter[28] ),
    .X(_300_));
 sky130_fd_sc_hd__and3b_2 _650_ (.A_N(_299_),
    .B(_300_),
    .C(_243_),
    .X(_020_));
 sky130_fd_sc_hd__or2_2 _651_ (.A(\counter[29] ),
    .B(_299_),
    .X(_301_));
 sky130_fd_sc_hd__nand2_2 _652_ (.A(\counter[29] ),
    .B(_299_),
    .Y(_302_));
 sky130_fd_sc_hd__and3_2 _653_ (.A(_243_),
    .B(_301_),
    .C(_302_),
    .X(_021_));
 sky130_fd_sc_hd__nand2_2 _654_ (.A(_092_),
    .B(_302_),
    .Y(_303_));
 sky130_fd_sc_hd__nor2_2 _655_ (.A(_092_),
    .B(_302_),
    .Y(_304_));
 sky130_fd_sc_hd__and3b_2 _656_ (.A_N(_304_),
    .B(_243_),
    .C(_303_),
    .X(_023_));
 sky130_fd_sc_hd__o21a_2 _657_ (.A1(\counter[31] ),
    .A2(_304_),
    .B1(_243_),
    .X(_024_));
 sky130_fd_sc_hd__and2_2 _658_ (.A(_078_),
    .B(\counter[28] ),
    .X(_305_));
 sky130_fd_sc_hd__and2_2 _659_ (.A(_090_),
    .B(\counter[29] ),
    .X(_306_));
 sky130_fd_sc_hd__a21oi_2 _660_ (.A1(_091_),
    .A2(\counter[30] ),
    .B1(\counter[31] ),
    .Y(_307_));
 sky130_fd_sc_hd__o22a_2 _661_ (.A1(_090_),
    .A2(\counter[29] ),
    .B1(\counter[28] ),
    .B2(_078_),
    .X(_308_));
 sky130_fd_sc_hd__o221a_2 _662_ (.A1(_091_),
    .A2(\counter[30] ),
    .B1(_093_),
    .B2(psc[28]),
    .C1(_307_),
    .X(_309_));
 sky130_fd_sc_hd__and4bb_2 _663_ (.A_N(_305_),
    .B_N(_306_),
    .C(_308_),
    .D(_309_),
    .X(_310_));
 sky130_fd_sc_hd__a22o_2 _664_ (.A1(psc[28]),
    .A2(_093_),
    .B1(_094_),
    .B2(psc[27]),
    .X(_311_));
 sky130_fd_sc_hd__a21oi_2 _665_ (.A1(_081_),
    .A2(\counter[24] ),
    .B1(_311_),
    .Y(_312_));
 sky130_fd_sc_hd__o22a_2 _666_ (.A1(_080_),
    .A2(\counter[25] ),
    .B1(\counter[24] ),
    .B2(_081_),
    .X(_313_));
 sky130_fd_sc_hd__a2bb2o_2 _667_ (.A1_N(psc[27]),
    .A2_N(_094_),
    .B1(\counter[25] ),
    .B2(_080_),
    .X(_314_));
 sky130_fd_sc_hd__inv_2 _668_ (.A(_314_),
    .Y(_315_));
 sky130_fd_sc_hd__and4_2 _669_ (.A(_310_),
    .B(_312_),
    .C(_313_),
    .D(_315_),
    .X(_316_));
 sky130_fd_sc_hd__and2_2 _670_ (.A(_082_),
    .B(\counter[23] ),
    .X(_317_));
 sky130_fd_sc_hd__nor2_2 _671_ (.A(_082_),
    .B(\counter[23] ),
    .Y(_318_));
 sky130_fd_sc_hd__or2_2 _672_ (.A(_083_),
    .B(\counter[22] ),
    .X(_319_));
 sky130_fd_sc_hd__and2_2 _673_ (.A(_083_),
    .B(\counter[22] ),
    .X(_320_));
 sky130_fd_sc_hd__a22o_2 _674_ (.A1(_084_),
    .A2(\counter[21] ),
    .B1(\counter[20] ),
    .B2(_085_),
    .X(_321_));
 sky130_fd_sc_hd__and2b_2 _675_ (.A_N(psc[20]),
    .B(\counter[19] ),
    .X(_322_));
 sky130_fd_sc_hd__nor2_2 _676_ (.A(_086_),
    .B(\counter[18] ),
    .Y(_323_));
 sky130_fd_sc_hd__nand2b_2 _677_ (.A_N(\counter[19] ),
    .B(psc[20]),
    .Y(_324_));
 sky130_fd_sc_hd__a21bo_2 _678_ (.A1(_086_),
    .A2(\counter[18] ),
    .B1_N(_324_),
    .X(_325_));
 sky130_fd_sc_hd__o22a_2 _679_ (.A1(_087_),
    .A2(\counter[17] ),
    .B1(\counter[16] ),
    .B2(_088_),
    .X(_326_));
 sky130_fd_sc_hd__and2_2 _680_ (.A(_087_),
    .B(\counter[17] ),
    .X(_327_));
 sky130_fd_sc_hd__o32a_2 _681_ (.A1(_325_),
    .A2(_326_),
    .A3(_327_),
    .B1(\counter[18] ),
    .B2(_086_),
    .X(_328_));
 sky130_fd_sc_hd__o221a_2 _682_ (.A1(_085_),
    .A2(\counter[20] ),
    .B1(_322_),
    .B2(_328_),
    .C1(_324_),
    .X(_329_));
 sky130_fd_sc_hd__o22a_2 _683_ (.A1(_084_),
    .A2(\counter[21] ),
    .B1(_321_),
    .B2(_329_),
    .X(_330_));
 sky130_fd_sc_hd__o221a_2 _684_ (.A1(_082_),
    .A2(\counter[23] ),
    .B1(_320_),
    .B2(_330_),
    .C1(_319_),
    .X(_331_));
 sky130_fd_sc_hd__nor2_2 _685_ (.A(_317_),
    .B(_331_),
    .Y(_332_));
 sky130_fd_sc_hd__or3b_2 _686_ (.A(_318_),
    .B(_321_),
    .C_N(_319_),
    .X(_333_));
 sky130_fd_sc_hd__nand2b_2 _687_ (.A_N(_325_),
    .B(_326_),
    .Y(_334_));
 sky130_fd_sc_hd__a2111o_2 _688_ (.A1(_088_),
    .A2(\counter[16] ),
    .B1(_322_),
    .C1(_323_),
    .D1(_327_),
    .X(_335_));
 sky130_fd_sc_hd__o22a_2 _689_ (.A1(_084_),
    .A2(\counter[21] ),
    .B1(\counter[20] ),
    .B2(_085_),
    .X(_336_));
 sky130_fd_sc_hd__or4b_2 _690_ (.A(_317_),
    .B(_320_),
    .C(_335_),
    .D_N(_336_),
    .X(_337_));
 sky130_fd_sc_hd__nor3_2 _691_ (.A(_333_),
    .B(_334_),
    .C(_337_),
    .Y(_338_));
 sky130_fd_sc_hd__nand2b_2 _692_ (.A_N(\counter[7] ),
    .B(psc[8]),
    .Y(_339_));
 sky130_fd_sc_hd__and2_2 _693_ (.A(_071_),
    .B(\counter[6] ),
    .X(_340_));
 sky130_fd_sc_hd__a22o_2 _694_ (.A1(_070_),
    .A2(\counter[5] ),
    .B1(\counter[4] ),
    .B2(_069_),
    .X(_341_));
 sky130_fd_sc_hd__and2b_2 _695_ (.A_N(psc[4]),
    .B(\counter[3] ),
    .X(_342_));
 sky130_fd_sc_hd__and2b_2 _696_ (.A_N(\counter[3] ),
    .B(psc[4]),
    .X(_343_));
 sky130_fd_sc_hd__xor2_2 _697_ (.A(psc[3]),
    .B(\counter[2] ),
    .X(_344_));
 sky130_fd_sc_hd__or3_2 _698_ (.A(_342_),
    .B(_343_),
    .C(_344_),
    .X(_345_));
 sky130_fd_sc_hd__nand2_2 _699_ (.A(_067_),
    .B(psc[2]),
    .Y(_346_));
 sky130_fd_sc_hd__a2bb2o_2 _700_ (.A1_N(_066_),
    .A2_N(psc[1]),
    .B1(\counter[1] ),
    .B2(_068_),
    .X(_347_));
 sky130_fd_sc_hd__a21o_2 _701_ (.A1(_346_),
    .A2(_347_),
    .B1(_345_),
    .X(_348_));
 sky130_fd_sc_hd__or3b_2 _702_ (.A(\counter[2] ),
    .B(_342_),
    .C_N(psc[3]),
    .X(_349_));
 sky130_fd_sc_hd__nor2_2 _703_ (.A(_069_),
    .B(\counter[4] ),
    .Y(_350_));
 sky130_fd_sc_hd__nor2_2 _704_ (.A(_343_),
    .B(_350_),
    .Y(_351_));
 sky130_fd_sc_hd__a31o_2 _705_ (.A1(_348_),
    .A2(_349_),
    .A3(_351_),
    .B1(_341_),
    .X(_352_));
 sky130_fd_sc_hd__o221a_2 _706_ (.A1(_071_),
    .A2(\counter[6] ),
    .B1(\counter[5] ),
    .B2(_070_),
    .C1(_352_),
    .X(_353_));
 sky130_fd_sc_hd__o21ai_2 _707_ (.A1(_340_),
    .A2(_353_),
    .B1(_339_),
    .Y(_354_));
 sky130_fd_sc_hd__a2bb2o_2 _708_ (.A1_N(\counter[8] ),
    .A2_N(_072_),
    .B1(psc[10]),
    .B2(_077_),
    .X(_355_));
 sky130_fd_sc_hd__o22a_2 _709_ (.A1(psc[14]),
    .A2(_074_),
    .B1(_075_),
    .B2(psc[13]),
    .X(_356_));
 sky130_fd_sc_hd__inv_2 _710_ (.A(_356_),
    .Y(_357_));
 sky130_fd_sc_hd__and2_2 _711_ (.A(psc[13]),
    .B(_075_),
    .X(_358_));
 sky130_fd_sc_hd__nand2b_2 _712_ (.A_N(\counter[11] ),
    .B(psc[12]),
    .Y(_359_));
 sky130_fd_sc_hd__o221a_2 _713_ (.A1(psc[11]),
    .A2(_076_),
    .B1(_077_),
    .B2(psc[10]),
    .C1(_359_),
    .X(_360_));
 sky130_fd_sc_hd__and2b_2 _714_ (.A_N(psc[12]),
    .B(\counter[11] ),
    .X(_361_));
 sky130_fd_sc_hd__nor2_2 _715_ (.A(\counter[15] ),
    .B(_089_),
    .Y(_362_));
 sky130_fd_sc_hd__o2bb2a_2 _716_ (.A1_N(\counter[15] ),
    .A2_N(_089_),
    .B1(_073_),
    .B2(psc[15]),
    .X(_363_));
 sky130_fd_sc_hd__a22o_2 _717_ (.A1(psc[15]),
    .A2(_073_),
    .B1(_074_),
    .B2(psc[14]),
    .X(_364_));
 sky130_fd_sc_hd__a221o_2 _718_ (.A1(psc[11]),
    .A2(_076_),
    .B1(\counter[8] ),
    .B2(_072_),
    .C1(_358_),
    .X(_365_));
 sky130_fd_sc_hd__nand2_2 _719_ (.A(_360_),
    .B(_363_),
    .Y(_366_));
 sky130_fd_sc_hd__or4_2 _720_ (.A(_355_),
    .B(_357_),
    .C(_364_),
    .D(_366_),
    .X(_367_));
 sky130_fd_sc_hd__or4_2 _721_ (.A(_361_),
    .B(_362_),
    .C(_365_),
    .D(_367_),
    .X(_368_));
 sky130_fd_sc_hd__nand2b_2 _722_ (.A_N(psc[8]),
    .B(\counter[7] ),
    .Y(_369_));
 sky130_fd_sc_hd__and3b_2 _723_ (.A_N(_368_),
    .B(_369_),
    .C(_354_),
    .X(_370_));
 sky130_fd_sc_hd__nand2b_2 _724_ (.A_N(_358_),
    .B(_361_),
    .Y(_371_));
 sky130_fd_sc_hd__a221o_2 _725_ (.A1(psc[11]),
    .A2(_076_),
    .B1(_355_),
    .B2(_360_),
    .C1(_358_),
    .X(_372_));
 sky130_fd_sc_hd__nand2_2 _726_ (.A(_371_),
    .B(_372_),
    .Y(_373_));
 sky130_fd_sc_hd__a21oi_2 _727_ (.A1(_359_),
    .A2(_373_),
    .B1(_357_),
    .Y(_374_));
 sky130_fd_sc_hd__o21a_2 _728_ (.A1(_364_),
    .A2(_374_),
    .B1(_363_),
    .X(_375_));
 sky130_fd_sc_hd__o31a_2 _729_ (.A1(_362_),
    .A2(_370_),
    .A3(_375_),
    .B1(_338_),
    .X(_376_));
 sky130_fd_sc_hd__o21a_2 _730_ (.A1(_332_),
    .A2(_376_),
    .B1(_316_),
    .X(_377_));
 sky130_fd_sc_hd__o21bai_2 _731_ (.A1(_313_),
    .A2(_314_),
    .B1_N(_311_),
    .Y(_378_));
 sky130_fd_sc_hd__o22ai_2 _732_ (.A1(_091_),
    .A2(\counter[30] ),
    .B1(_306_),
    .B2(_308_),
    .Y(_379_));
 sky130_fd_sc_hd__a22o_2 _733_ (.A1(_310_),
    .A2(_378_),
    .B1(_379_),
    .B2(_307_),
    .X(_380_));
 sky130_fd_sc_hd__o221a_2 _734_ (.A1(_071_),
    .A2(\counter[6] ),
    .B1(\counter[5] ),
    .B2(_070_),
    .C1(_369_),
    .X(_381_));
 sky130_fd_sc_hd__or4bb_2 _735_ (.A(_341_),
    .B(_347_),
    .C_N(_381_),
    .D_N(_339_),
    .X(_382_));
 sky130_fd_sc_hd__a2111o_2 _736_ (.A1(_066_),
    .A2(psc[1]),
    .B1(_340_),
    .C1(_345_),
    .D1(_350_),
    .X(_383_));
 sky130_fd_sc_hd__or3b_2 _737_ (.A(_382_),
    .B(_383_),
    .C_N(_346_),
    .X(_384_));
 sky130_fd_sc_hd__nand2_2 _738_ (.A(_316_),
    .B(_338_),
    .Y(_385_));
 sky130_fd_sc_hd__o32a_2 _739_ (.A1(_368_),
    .A2(_384_),
    .A3(_385_),
    .B1(_377_),
    .B2(_380_),
    .X(_032_));
 sky130_fd_sc_hd__inv_2 _740_ (.A(rst),
    .Y(_034_));
 sky130_fd_sc_hd__inv_2 _741_ (.A(rst),
    .Y(_035_));
 sky130_fd_sc_hd__inv_2 _742_ (.A(rst),
    .Y(_036_));
 sky130_fd_sc_hd__inv_2 _743_ (.A(rst),
    .Y(_037_));
 sky130_fd_sc_hd__inv_2 _744_ (.A(rst),
    .Y(_038_));
 sky130_fd_sc_hd__inv_2 _745_ (.A(rst),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _746_ (.A(rst),
    .Y(_040_));
 sky130_fd_sc_hd__inv_2 _747_ (.A(rst),
    .Y(_041_));
 sky130_fd_sc_hd__inv_2 _748_ (.A(rst),
    .Y(_042_));
 sky130_fd_sc_hd__inv_2 _749_ (.A(rst),
    .Y(_043_));
 sky130_fd_sc_hd__inv_2 _750_ (.A(rst),
    .Y(_044_));
 sky130_fd_sc_hd__inv_2 _751_ (.A(rst),
    .Y(_045_));
 sky130_fd_sc_hd__inv_2 _752_ (.A(rst),
    .Y(_046_));
 sky130_fd_sc_hd__inv_2 _753_ (.A(rst),
    .Y(_047_));
 sky130_fd_sc_hd__inv_2 _754_ (.A(rst),
    .Y(_048_));
 sky130_fd_sc_hd__inv_2 _755_ (.A(rst),
    .Y(_049_));
 sky130_fd_sc_hd__inv_2 _756_ (.A(rst),
    .Y(_050_));
 sky130_fd_sc_hd__inv_2 _757_ (.A(rst),
    .Y(_051_));
 sky130_fd_sc_hd__inv_2 _758_ (.A(rst),
    .Y(_052_));
 sky130_fd_sc_hd__inv_2 _759_ (.A(rst),
    .Y(_053_));
 sky130_fd_sc_hd__inv_2 _760_ (.A(rst),
    .Y(_054_));
 sky130_fd_sc_hd__inv_2 _761_ (.A(rst),
    .Y(_055_));
 sky130_fd_sc_hd__inv_2 _762_ (.A(rst),
    .Y(_056_));
 sky130_fd_sc_hd__inv_2 _763_ (.A(rst),
    .Y(_057_));
 sky130_fd_sc_hd__inv_2 _764_ (.A(rst),
    .Y(_058_));
 sky130_fd_sc_hd__inv_2 _765_ (.A(rst),
    .Y(_059_));
 sky130_fd_sc_hd__inv_2 _766_ (.A(rst),
    .Y(_060_));
 sky130_fd_sc_hd__inv_2 _767_ (.A(rst),
    .Y(_061_));
 sky130_fd_sc_hd__inv_2 _768_ (.A(rst),
    .Y(_062_));
 sky130_fd_sc_hd__inv_2 _769_ (.A(rst),
    .Y(_063_));
 sky130_fd_sc_hd__inv_2 _770_ (.A(rst),
    .Y(_064_));
 sky130_fd_sc_hd__inv_2 _771_ (.A(rst),
    .Y(_065_));
 sky130_fd_sc_hd__dfrtp_2 _772_ (.CLK(clk),
    .D(_032_),
    .RESET_B(_033_),
    .Q(out));
 sky130_fd_sc_hd__dfrtp_2 _773_ (.CLK(clk),
    .D(_000_),
    .RESET_B(_034_),
    .Q(\counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _774_ (.CLK(clk),
    .D(_011_),
    .RESET_B(_035_),
    .Q(\counter[1] ));
 sky130_fd_sc_hd__dfrtp_2 _775_ (.CLK(clk),
    .D(_022_),
    .RESET_B(_036_),
    .Q(\counter[2] ));
 sky130_fd_sc_hd__dfrtp_2 _776_ (.CLK(clk),
    .D(_025_),
    .RESET_B(_037_),
    .Q(\counter[3] ));
 sky130_fd_sc_hd__dfrtp_2 _777_ (.CLK(clk),
    .D(_026_),
    .RESET_B(_038_),
    .Q(\counter[4] ));
 sky130_fd_sc_hd__dfrtp_2 _778_ (.CLK(clk),
    .D(_027_),
    .RESET_B(_039_),
    .Q(\counter[5] ));
 sky130_fd_sc_hd__dfrtp_2 _779_ (.CLK(clk),
    .D(_028_),
    .RESET_B(_040_),
    .Q(\counter[6] ));
 sky130_fd_sc_hd__dfrtp_2 _780_ (.CLK(clk),
    .D(_029_),
    .RESET_B(_041_),
    .Q(\counter[7] ));
 sky130_fd_sc_hd__dfrtp_2 _781_ (.CLK(clk),
    .D(_030_),
    .RESET_B(_042_),
    .Q(\counter[8] ));
 sky130_fd_sc_hd__dfrtp_2 _782_ (.CLK(clk),
    .D(_031_),
    .RESET_B(_043_),
    .Q(\counter[9] ));
 sky130_fd_sc_hd__dfrtp_2 _783_ (.CLK(clk),
    .D(_001_),
    .RESET_B(_044_),
    .Q(\counter[10] ));
 sky130_fd_sc_hd__dfrtp_2 _784_ (.CLK(clk),
    .D(_002_),
    .RESET_B(_045_),
    .Q(\counter[11] ));
 sky130_fd_sc_hd__dfrtp_2 _785_ (.CLK(clk),
    .D(_003_),
    .RESET_B(_046_),
    .Q(\counter[12] ));
 sky130_fd_sc_hd__dfrtp_2 _786_ (.CLK(clk),
    .D(_004_),
    .RESET_B(_047_),
    .Q(\counter[13] ));
 sky130_fd_sc_hd__dfrtp_2 _787_ (.CLK(clk),
    .D(_005_),
    .RESET_B(_048_),
    .Q(\counter[14] ));
 sky130_fd_sc_hd__dfrtp_2 _788_ (.CLK(clk),
    .D(_006_),
    .RESET_B(_049_),
    .Q(\counter[15] ));
 sky130_fd_sc_hd__dfrtp_2 _789_ (.CLK(clk),
    .D(_007_),
    .RESET_B(_050_),
    .Q(\counter[16] ));
 sky130_fd_sc_hd__dfrtp_2 _790_ (.CLK(clk),
    .D(_008_),
    .RESET_B(_051_),
    .Q(\counter[17] ));
 sky130_fd_sc_hd__dfrtp_2 _791_ (.CLK(clk),
    .D(_009_),
    .RESET_B(_052_),
    .Q(\counter[18] ));
 sky130_fd_sc_hd__dfrtp_2 _792_ (.CLK(clk),
    .D(_010_),
    .RESET_B(_053_),
    .Q(\counter[19] ));
 sky130_fd_sc_hd__dfrtp_2 _793_ (.CLK(clk),
    .D(_012_),
    .RESET_B(_054_),
    .Q(\counter[20] ));
 sky130_fd_sc_hd__dfrtp_2 _794_ (.CLK(clk),
    .D(_013_),
    .RESET_B(_055_),
    .Q(\counter[21] ));
 sky130_fd_sc_hd__dfrtp_2 _795_ (.CLK(clk),
    .D(_014_),
    .RESET_B(_056_),
    .Q(\counter[22] ));
 sky130_fd_sc_hd__dfrtp_2 _796_ (.CLK(clk),
    .D(_015_),
    .RESET_B(_057_),
    .Q(\counter[23] ));
 sky130_fd_sc_hd__dfrtp_2 _797_ (.CLK(clk),
    .D(_016_),
    .RESET_B(_058_),
    .Q(\counter[24] ));
 sky130_fd_sc_hd__dfrtp_2 _798_ (.CLK(clk),
    .D(_017_),
    .RESET_B(_059_),
    .Q(\counter[25] ));
 sky130_fd_sc_hd__dfrtp_2 _799_ (.CLK(clk),
    .D(_018_),
    .RESET_B(_060_),
    .Q(\counter[26] ));
 sky130_fd_sc_hd__dfrtp_2 _800_ (.CLK(clk),
    .D(_019_),
    .RESET_B(_061_),
    .Q(\counter[27] ));
 sky130_fd_sc_hd__dfrtp_2 _801_ (.CLK(clk),
    .D(_020_),
    .RESET_B(_062_),
    .Q(\counter[28] ));
 sky130_fd_sc_hd__dfrtp_2 _802_ (.CLK(clk),
    .D(_021_),
    .RESET_B(_063_),
    .Q(\counter[29] ));
 sky130_fd_sc_hd__dfrtp_2 _803_ (.CLK(clk),
    .D(_023_),
    .RESET_B(_064_),
    .Q(\counter[30] ));
 sky130_fd_sc_hd__dfrtp_2 _804_ (.CLK(clk),
    .D(_024_),
    .RESET_B(_065_),
    .Q(\counter[31] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_165 ();
endmodule
