VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO freq_psc
  CLASS BLOCK ;
  FOREIGN freq_psc ;
  ORIGIN 0.000 0.000 ;
  SIZE 72.390 BY 83.110 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 70.960 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 70.960 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END clk
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END out
  PIN psc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 68.390 47.640 72.390 48.240 ;
    END
  END psc[0]
  PIN psc[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 79.110 26.130 83.110 ;
    END
  END psc[10]
  PIN psc[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 79.110 29.350 83.110 ;
    END
  END psc[11]
  PIN psc[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END psc[12]
  PIN psc[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END psc[13]
  PIN psc[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END psc[14]
  PIN psc[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END psc[15]
  PIN psc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 68.390 51.040 72.390 51.640 ;
    END
  END psc[1]
  PIN psc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 68.390 44.240 72.390 44.840 ;
    END
  END psc[2]
  PIN psc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 68.390 54.440 72.390 55.040 ;
    END
  END psc[3]
  PIN psc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 79.110 48.670 83.110 ;
    END
  END psc[4]
  PIN psc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 79.110 45.450 83.110 ;
    END
  END psc[5]
  PIN psc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 38.730 79.110 39.010 83.110 ;
    END
  END psc[6]
  PIN psc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 79.110 35.790 83.110 ;
    END
  END psc[7]
  PIN psc[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 79.110 42.230 83.110 ;
    END
  END psc[8]
  PIN psc[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 79.110 32.570 83.110 ;
    END
  END psc[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 68.390 17.040 72.390 17.640 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 66.890 70.805 ;
      LAYER li1 ;
        RECT 5.520 10.795 66.700 70.805 ;
      LAYER met1 ;
        RECT 4.210 10.640 66.700 70.960 ;
      LAYER met2 ;
        RECT 4.230 78.830 25.570 79.110 ;
        RECT 26.410 78.830 28.790 79.110 ;
        RECT 29.630 78.830 32.010 79.110 ;
        RECT 32.850 78.830 35.230 79.110 ;
        RECT 36.070 78.830 38.450 79.110 ;
        RECT 39.290 78.830 41.670 79.110 ;
        RECT 42.510 78.830 44.890 79.110 ;
        RECT 45.730 78.830 48.110 79.110 ;
        RECT 48.950 78.830 65.230 79.110 ;
        RECT 4.230 4.280 65.230 78.830 ;
        RECT 4.230 4.000 25.570 4.280 ;
        RECT 26.410 4.000 28.790 4.280 ;
        RECT 29.630 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 65.230 4.280 ;
      LAYER met3 ;
        RECT 3.990 55.440 68.390 70.885 ;
        RECT 3.990 54.040 67.990 55.440 ;
        RECT 3.990 52.040 68.390 54.040 ;
        RECT 3.990 50.640 67.990 52.040 ;
        RECT 3.990 48.640 68.390 50.640 ;
        RECT 4.400 47.240 67.990 48.640 ;
        RECT 3.990 45.240 68.390 47.240 ;
        RECT 3.990 43.840 67.990 45.240 ;
        RECT 3.990 31.640 68.390 43.840 ;
        RECT 4.400 30.240 68.390 31.640 ;
        RECT 3.990 18.040 68.390 30.240 ;
        RECT 3.990 16.640 67.990 18.040 ;
        RECT 3.990 10.715 68.390 16.640 ;
  END
END freq_psc
END LIBRARY

