magic
tech sky130A
magscale 1 2
timestamp 1730308856
<< nwell >>
rect 1762 782 1968 1103
rect 594 1 848 491
rect 1792 260 1968 782
rect 594 0 835 1
rect 1429 -306 1432 260
rect 1765 -1 1968 260
rect 1792 -306 1968 -1
<< viali >>
rect 1507 736 1542 771
rect 1694 725 1728 759
rect 1509 272 1543 306
rect 1694 282 1728 316
rect 1489 -357 1534 -312
rect 1679 -351 1719 -311
rect 1821 -352 1861 -312
<< metal1 >>
rect 71 1162 124 1168
rect 1464 1109 1470 1162
rect 1523 1113 1529 1162
rect 1523 1109 1901 1113
rect 71 829 124 1109
rect 584 1069 656 1096
rect 584 1016 594 1069
rect 646 1016 656 1069
rect 1470 1060 1901 1109
rect 1681 1017 1901 1060
rect 1954 1017 1964 1113
rect 1395 771 1554 777
rect 1395 736 1507 771
rect 1542 736 1554 771
rect 1815 768 1867 774
rect 1395 730 1554 736
rect 1682 759 1815 765
rect 1395 548 1442 730
rect 1682 725 1694 759
rect 1728 725 1815 759
rect 1682 719 1815 725
rect 1815 710 1867 716
rect 1109 501 1442 548
rect 1489 494 1499 546
rect 1551 494 1561 546
rect 1732 325 1784 331
rect 1682 316 1732 322
rect 1299 306 1555 312
rect 1299 272 1509 306
rect 1543 272 1555 306
rect 1682 282 1694 316
rect 1728 282 1732 316
rect 1682 276 1732 282
rect 1299 266 1555 272
rect 1732 267 1784 273
rect 1225 -71 1484 -25
rect 1891 -71 1901 25
rect 1954 -71 1964 25
rect 1673 -305 1725 -299
rect 1477 -363 1483 -306
rect 1540 -363 1546 -306
rect 1673 -363 1725 -357
rect 1809 -358 1815 -306
rect 1867 -358 1873 -306
rect 773 -578 783 -525
rect 835 -578 845 -525
rect 773 -606 845 -578
rect 1470 -600 1535 -598
rect 1474 -601 1539 -600
rect 1470 -618 1543 -601
rect 1470 -671 1480 -618
rect 1533 -671 1543 -618
<< via1 >>
rect 71 1109 124 1162
rect 1470 1109 1523 1162
rect 594 1016 646 1069
rect 1901 1017 1954 1113
rect 1815 716 1867 768
rect 1499 494 1551 546
rect 1732 273 1784 325
rect 1901 -71 1954 25
rect 1483 -312 1540 -306
rect 1483 -357 1489 -312
rect 1489 -357 1534 -312
rect 1534 -357 1540 -312
rect 1483 -363 1540 -357
rect 1673 -311 1725 -305
rect 1673 -351 1679 -311
rect 1679 -351 1719 -311
rect 1719 -351 1725 -311
rect 1673 -357 1725 -351
rect 1815 -312 1867 -306
rect 1815 -352 1821 -312
rect 1821 -352 1861 -312
rect 1861 -352 1867 -312
rect 1815 -358 1867 -352
rect 783 -578 835 -525
rect 1480 -671 1533 -618
<< metal2 >>
rect 1470 1162 1523 1168
rect 65 1109 71 1162
rect 124 1109 1470 1162
rect 1470 1103 1523 1109
rect 1901 1113 1954 1123
rect 592 1071 648 1081
rect 592 1004 648 1014
rect 690 932 722 953
rect 1007 546 1059 805
rect 1809 716 1815 768
rect 1867 716 1873 768
rect 1499 546 1551 556
rect 1007 494 1499 546
rect 1007 434 1059 494
rect 1499 484 1551 494
rect 682 382 1059 434
rect 682 66 734 382
rect 1726 273 1732 325
rect 1784 273 1790 325
rect 377 14 734 66
rect 377 -314 429 14
rect 1483 -306 1540 -300
rect 1735 -305 1781 273
rect 1818 -300 1864 716
rect 1901 25 1954 1017
rect 1901 -81 1954 -71
rect 1366 -363 1483 -306
rect 1667 -357 1673 -305
rect 1725 -354 1781 -305
rect 1815 -306 1867 -300
rect 1725 -357 1731 -354
rect 429 -618 482 -405
rect 718 -474 756 -449
rect 781 -523 837 -513
rect 1366 -523 1423 -363
rect 1483 -369 1540 -363
rect 1815 -364 1867 -358
rect 837 -580 1423 -523
rect 781 -590 837 -580
rect 1480 -618 1533 -608
rect 429 -671 1480 -618
rect 1480 -681 1533 -671
<< via2 >>
rect 592 1069 648 1071
rect 592 1016 594 1069
rect 594 1016 646 1069
rect 646 1016 648 1069
rect 592 1014 648 1016
rect 781 -525 837 -523
rect 781 -578 783 -525
rect 783 -578 835 -525
rect 835 -578 837 -525
rect 781 -580 837 -578
<< metal3 >>
rect 582 1071 658 1076
rect 582 1014 592 1071
rect 648 1014 658 1071
rect 582 1009 658 1014
rect 590 276 650 1009
rect 590 215 839 276
rect 779 -518 839 215
rect 771 -523 847 -518
rect 771 -580 781 -523
rect 837 -580 847 -523
rect 771 -585 847 -580
use tspc_dff  x1
timestamp 1730306127
transform 1 0 697 0 1 60
box -697 -60 635 1065
use tspc_dff  x2
timestamp 1730306127
transform -1 0 732 0 -1 431
box -697 -60 635 1065
use sky130_fd_sc_hd__and2_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform -1 0 1930 0 1 -567
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730246015
transform 1 0 1470 0 -1 521
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x5
timestamp 1730246015
transform 1 0 1470 0 1 521
box -38 -48 314 592
<< labels >>
flabel metal2 1147 -651 1147 -651 0 FreeSans 160 0 0 0 DVSS
port 0 nsew
flabel metal2 1925 607 1925 607 0 FreeSans 160 90 0 0 DVDD
port 1 nsew
flabel metal2 1837 -228 1837 -228 0 FreeSans 160 0 0 0 U
port 2 nsew
flabel metal2 1758 -266 1758 -266 0 FreeSans 160 0 0 0 D
port 3 nsew
flabel metal2 707 943 707 943 0 FreeSans 160 0 0 0 vin1
port 4 nsew
flabel metal2 741 -461 741 -461 0 FreeSans 160 0 0 0 vin2
port 5 nsew
<< end >>
