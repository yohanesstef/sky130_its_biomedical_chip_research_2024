magic
tech sky130A
magscale 1 2
timestamp 1730039636
<< nwell >>
rect 2703 2534 3590 2855
rect 2418 1446 2439 2012
<< nsubdiff >>
rect 3472 2716 3554 2740
rect 3472 2682 3496 2716
rect 3530 2682 3554 2716
rect 3472 2658 3554 2682
<< nsubdiffcont >>
rect 3496 2682 3530 2716
<< locali >>
rect 3472 2716 3554 2740
rect 3472 2682 3496 2716
rect 3530 2682 3554 2716
rect 3472 2658 3554 2682
rect 2973 2470 3066 2544
<< viali >>
rect 3496 2682 3530 2716
rect 2759 2491 2793 2525
rect 3228 2488 3262 2522
rect 3358 2488 3392 2522
rect 2503 2019 2703 2057
rect 3332 2023 3366 2057
rect 2492 1403 2712 1437
rect 3328 1397 3368 1437
<< metal1 >>
rect 933 2824 1408 2875
rect 2164 2829 2625 2875
rect 933 1167 984 2824
rect 1043 2397 1053 2625
rect 1105 2397 1115 2625
rect 2195 2503 2517 2555
rect 2092 2250 2437 2299
rect 2465 2274 2517 2503
rect 2579 2531 2625 2829
rect 2760 2791 2770 2843
rect 2988 2791 2998 2843
rect 3459 2769 3767 2865
rect 3484 2716 3542 2769
rect 3484 2682 3496 2716
rect 3530 2682 3542 2716
rect 3484 2676 3542 2682
rect 2579 2525 2805 2531
rect 2579 2491 2759 2525
rect 2793 2491 2805 2525
rect 2579 2485 2805 2491
rect 3209 2479 3219 2531
rect 3271 2479 3281 2531
rect 3346 2522 3643 2528
rect 3346 2488 3358 2522
rect 3392 2488 3643 2522
rect 3346 2482 3643 2488
rect 2294 2040 2340 2067
rect 2388 2063 2437 2250
rect 3487 2247 3497 2299
rect 3549 2247 3559 2299
rect 3597 2063 3643 2482
rect 2388 2057 2715 2063
rect 2281 1812 2291 2040
rect 2343 1812 2353 2040
rect 2388 2019 2503 2057
rect 2703 2019 2715 2057
rect 2388 2014 2715 2019
rect 3320 2057 3643 2063
rect 3320 2023 3332 2057
rect 3366 2023 3643 2057
rect 3320 2017 3643 2023
rect 2491 2013 2715 2014
rect 3671 1777 3767 2769
rect 2322 1725 2711 1777
rect 2288 1681 2711 1725
rect 3535 1681 3767 1777
rect 2288 1602 2418 1681
rect 2322 1583 2418 1602
rect 2482 1443 2492 1446
rect 2480 1397 2492 1443
rect 2712 1443 2722 1446
rect 2482 1394 2492 1397
rect 2712 1397 2724 1443
rect 2712 1394 2722 1397
rect 3316 1391 3322 1443
rect 3374 1391 3380 1443
rect 933 1116 1273 1167
rect 2484 1159 2494 1211
rect 2712 1159 2722 1211
rect 3491 1159 3497 1211
rect 3549 1159 3555 1211
<< via1 >>
rect 1053 2397 1105 2625
rect 2770 2791 2988 2843
rect 3219 2522 3271 2531
rect 3219 2488 3228 2522
rect 3228 2488 3262 2522
rect 3262 2488 3271 2522
rect 3219 2479 3271 2488
rect 3497 2247 3549 2299
rect 2291 1812 2343 2040
rect 2492 1437 2712 1446
rect 2492 1403 2712 1437
rect 2492 1394 2712 1403
rect 3322 1437 3374 1443
rect 3322 1397 3328 1437
rect 3328 1397 3368 1437
rect 3368 1397 3374 1437
rect 3322 1391 3374 1397
rect 2494 1159 2712 1211
rect 3497 1159 3549 1211
<< metal2 >>
rect 1029 2843 3009 2865
rect 1029 2791 2770 2843
rect 2988 2791 3009 2843
rect 1029 2769 3009 2791
rect 1029 2625 1125 2769
rect 1583 2683 1600 2714
rect 1029 2397 1053 2625
rect 1105 2397 1125 2625
rect 3219 2531 3271 2541
rect 3271 2479 3469 2531
rect 3219 2469 3271 2479
rect 1029 2387 1125 2397
rect 2291 2040 2343 2050
rect 2343 1815 2475 1861
rect 2291 1802 2343 1812
rect 2429 1456 2475 1815
rect 2429 1446 2712 1456
rect 2429 1394 2492 1446
rect 3322 1443 3374 1449
rect 3417 1443 3469 2479
rect 2712 1397 2724 1443
rect 2429 1384 2712 1394
rect 3374 1391 3469 1443
rect 3497 2299 3549 2309
rect 3322 1385 3374 1391
rect 1424 1210 1477 1345
rect 1812 1290 1822 1302
rect 2494 1211 2712 1221
rect 1424 1159 2494 1210
rect 3497 1211 3549 2247
rect 2712 1159 2741 1210
rect 1424 1157 2741 1159
rect 2494 1149 2712 1157
rect 3497 1153 3549 1159
use tspc_dff  x1
timestamp 1730031749
transform 1 0 1679 0 1 1810
box -697 -60 635 1065
use tspc_dff  x2
timestamp 1730031749
transform -1 0 1727 0 -1 2181
box -697 -60 635 1065
use sky130_fd_sc_hd__and2_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3477 0 1 2273
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2465 0 -1 2273
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  x5
timestamp 1704896540
transform 1 0 2465 0 1 1185
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  x6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3017 0 1 2273
box -38 -48 314 592
<< labels >>
flabel metal1 3717 1772 3717 1772 0 FreeSans 1600 0 0 0 DVDD
port 0 nsew
flabel metal2 2106 1174 2106 1174 0 FreeSans 1600 0 0 0 DVSS
port 1 nsew
flabel metal2 3295 2505 3295 2505 0 FreeSans 1600 0 0 0 D
port 3 nsew
flabel metal2 1591 2697 1591 2697 0 FreeSans 1600 0 0 0 VIN1
port 4 nsew
flabel metal2 1816 1296 1816 1296 0 FreeSans 1600 0 0 0 VIN2
port 5 nsew
flabel metal1 3512 2498 3512 2498 0 FreeSans 1600 0 0 0 U
port 2 nsew
<< end >>
