magic
tech sky130A
timestamp 1730127321
<< nmos >>
rect -60 -500 60 500
<< ndiff >>
rect -89 494 -60 500
rect -89 -494 -83 494
rect -66 -494 -60 494
rect -89 -500 -60 -494
rect 60 494 89 500
rect 60 -494 66 494
rect 83 -494 89 494
rect 60 -500 89 -494
<< ndiffc >>
rect -83 -494 -66 494
rect 66 -494 83 494
<< poly >>
rect -60 536 60 544
rect -60 519 -52 536
rect 52 519 60 536
rect -60 500 60 519
rect -60 -519 60 -500
rect -60 -536 -52 -519
rect 52 -536 60 -519
rect -60 -544 60 -536
<< polycont >>
rect -52 519 52 536
rect -52 -536 52 -519
<< locali >>
rect -60 519 -52 536
rect 52 519 60 536
rect -83 494 -66 502
rect -83 -502 -66 -494
rect 66 494 83 502
rect 66 -502 83 -494
rect -60 -536 -52 -519
rect 52 -536 60 -519
<< viali >>
rect -52 519 52 536
rect -83 -494 -66 494
rect 66 -494 83 494
rect -52 -536 52 -519
<< metal1 >>
rect -58 536 58 539
rect -58 519 -52 536
rect 52 519 58 536
rect -58 516 58 519
rect -86 494 -63 500
rect -86 -494 -83 494
rect -66 -494 -63 494
rect -86 -500 -63 -494
rect 63 494 86 500
rect 63 -494 66 494
rect 83 -494 86 494
rect 63 -500 86 -494
rect -58 -519 58 -516
rect -58 -536 -52 -519
rect 52 -536 58 -519
rect -58 -539 58 -536
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
