magic
tech sky130A
magscale 1 2
timestamp 1729853601
<< nwell >>
rect -183 498 348 1211
rect -183 464 166 498
rect 178 464 348 498
rect -183 -127 348 464
<< nsubdiff >>
rect -147 1141 -87 1175
rect 252 1141 312 1175
rect -147 1115 -113 1141
rect 278 1115 312 1141
rect -147 -57 -113 -31
rect 278 -57 312 -31
rect -147 -91 -87 -57
rect 252 -91 312 -57
<< nsubdiffcont >>
rect -87 1141 252 1175
rect -147 -31 -113 1115
rect 278 -31 312 1115
rect -87 -91 252 -57
<< poly >>
rect -62 1103 36 1119
rect -62 1069 -46 1103
rect -12 1069 36 1103
rect -62 1053 36 1069
rect 0 1044 36 1053
<< polycont >>
rect -46 1069 -12 1103
<< locali >>
rect -147 1141 -87 1175
rect 252 1141 312 1175
rect -147 1115 -113 1141
rect 278 1115 312 1141
rect -62 1069 -46 1103
rect -12 1069 4 1103
rect -147 -57 -113 -31
rect 278 -57 312 -31
rect -147 -91 -87 -57
rect 252 -91 312 -57
<< viali >>
rect 48 1141 82 1175
rect -497 303 -463 337
rect -46 1069 -12 1103
rect 592 248 626 282
<< metal1 >>
rect 36 1175 94 1181
rect 36 1141 48 1175
rect 82 1141 94 1175
rect 36 1135 94 1141
rect -451 1103 4 1119
rect -451 1069 -46 1103
rect -12 1069 4 1103
rect -451 1053 4 1069
rect -451 639 -379 1053
rect 42 1010 88 1135
rect 529 628 595 681
rect -370 494 -12 528
rect 178 464 532 498
rect -503 343 -457 427
rect -509 337 -451 343
rect -509 303 -497 337
rect -463 303 -451 337
rect -509 297 -451 303
rect 586 288 632 372
rect 580 282 638 288
rect 580 248 592 282
rect 626 248 638 282
rect 580 242 638 248
rect -46 84 -12 112
rect -46 15 -12 74
rect -46 -19 162 15
use sky130_fd_pr__pfet_01v8_2V7TNJ  sky130_fd_pr__pfet_01v8_2V7TNJ_0
timestamp 1729851530
transform 1 0 18 0 1 542
box -112 -542 112 542
use sky130_fd_pr__pfet_01v8_77ASL4  sky130_fd_pr__pfet_01v8_77ASL4_0
timestamp 1729851530
transform 1 0 130 0 1 506
box -130 -544 130 578
use sky130_fd_pr__nfet_01v8_4N4BM2  XM2
timestamp 1729853601
transform 1 0 -415 0 1 542
box -232 -275 232 275
use sky130_fd_pr__nfet_01v8_R32FGG  XM4
timestamp 1729853601
transform 1 0 562 0 1 511
box -214 -299 214 299
<< labels >>
flabel metal1 -413 1070 -413 1070 0 FreeSans 1600 0 0 0 U
port 0 nsew
flabel metal1 537 655 537 655 0 FreeSans 160 0 0 0 D
port 2 nsew
flabel metal1 357 481 357 481 0 FreeSans 800 0 0 0 VCON
port 3 nsew
flabel metal1 66 1123 66 1123 0 FreeSans 800 0 0 0 VDD
port 4 nsew
flabel metal1 -484 365 -484 365 0 FreeSans 800 0 0 0 GND
port 5 nsew
<< end >>
