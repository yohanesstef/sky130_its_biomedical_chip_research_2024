magic
tech sky130A
magscale 1 2
timestamp 1730455722
<< viali >>
rect 9873 14569 9907 14603
rect 6745 14433 6779 14467
rect 6193 14365 6227 14399
rect 6469 14365 6503 14399
rect 7205 14365 7239 14399
rect 8493 14365 8527 14399
rect 10057 14365 10091 14399
rect 6009 14229 6043 14263
rect 7389 14229 7423 14263
rect 8677 14229 8711 14263
rect 9137 14025 9171 14059
rect 10333 14025 10367 14059
rect 6745 13957 6779 13991
rect 6377 13889 6411 13923
rect 6561 13889 6595 13923
rect 7021 13889 7055 13923
rect 8953 13889 8987 13923
rect 9505 13889 9539 13923
rect 9597 13889 9631 13923
rect 10149 13889 10183 13923
rect 5457 13821 5491 13855
rect 6837 13821 6871 13855
rect 9689 13821 9723 13855
rect 9965 13821 9999 13855
rect 5825 13753 5859 13787
rect 6377 13753 6411 13787
rect 5917 13685 5951 13719
rect 6745 13685 6779 13719
rect 7205 13685 7239 13719
rect 8861 13685 8895 13719
rect 5273 13481 5307 13515
rect 6266 13481 6300 13515
rect 8953 13481 8987 13515
rect 4905 13413 4939 13447
rect 6009 13345 6043 13379
rect 7757 13345 7791 13379
rect 10425 13345 10459 13379
rect 10701 13345 10735 13379
rect 1409 13277 1443 13311
rect 4077 13277 4111 13311
rect 4537 13277 4571 13311
rect 4721 13277 4755 13311
rect 4813 13277 4847 13311
rect 5089 13277 5123 13311
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 5733 13277 5767 13311
rect 7849 13277 7883 13311
rect 8033 13277 8067 13311
rect 8217 13277 8251 13311
rect 8401 13277 8435 13311
rect 8585 13277 8619 13311
rect 5641 13209 5675 13243
rect 1593 13141 1627 13175
rect 3893 13141 3927 13175
rect 4629 13141 4663 13175
rect 5917 13141 5951 13175
rect 8769 13141 8803 13175
rect 6009 12937 6043 12971
rect 8493 12937 8527 12971
rect 9781 12937 9815 12971
rect 13277 12937 13311 12971
rect 2605 12869 2639 12903
rect 5181 12869 5215 12903
rect 6653 12869 6687 12903
rect 7113 12869 7147 12903
rect 8033 12869 8067 12903
rect 4997 12801 5031 12835
rect 5273 12801 5307 12835
rect 5641 12801 5675 12835
rect 6837 12801 6871 12835
rect 8401 12801 8435 12835
rect 8585 12801 8619 12835
rect 8953 12801 8987 12835
rect 10149 12801 10183 12835
rect 2789 12733 2823 12767
rect 2881 12733 2915 12767
rect 3249 12733 3283 12767
rect 4813 12733 4847 12767
rect 5549 12733 5583 12767
rect 5733 12733 5767 12767
rect 5825 12733 5859 12767
rect 6561 12733 6595 12767
rect 7573 12733 7607 12767
rect 8677 12733 8711 12767
rect 10057 12733 10091 12767
rect 11529 12733 11563 12767
rect 11805 12733 11839 12767
rect 7665 12665 7699 12699
rect 9689 12665 9723 12699
rect 4675 12597 4709 12631
rect 7205 12597 7239 12631
rect 7113 12393 7147 12427
rect 9413 12393 9447 12427
rect 3525 12325 3559 12359
rect 7297 12325 7331 12359
rect 10609 12325 10643 12359
rect 1409 12257 1443 12291
rect 4813 12257 4847 12291
rect 5549 12257 5583 12291
rect 7021 12257 7055 12291
rect 10333 12257 10367 12291
rect 1777 12189 1811 12223
rect 3341 12189 3375 12223
rect 3525 12189 3559 12223
rect 3893 12189 3927 12223
rect 4077 12189 4111 12223
rect 5273 12189 5307 12223
rect 7665 12189 7699 12223
rect 7819 12189 7853 12223
rect 9321 12189 9355 12223
rect 9505 12189 9539 12223
rect 10241 12189 10275 12223
rect 7573 12121 7607 12155
rect 3203 12053 3237 12087
rect 8033 12053 8067 12087
rect 1501 11849 1535 11883
rect 2145 11849 2179 11883
rect 2605 11849 2639 11883
rect 7113 11849 7147 11883
rect 7389 11849 7423 11883
rect 10793 11849 10827 11883
rect 1685 11713 1719 11747
rect 1777 11713 1811 11747
rect 2513 11713 2547 11747
rect 3065 11713 3099 11747
rect 5733 11713 5767 11747
rect 5917 11713 5951 11747
rect 6377 11713 6411 11747
rect 6745 11713 6779 11747
rect 7665 11713 7699 11747
rect 7849 11713 7883 11747
rect 8769 11713 8803 11747
rect 2789 11645 2823 11679
rect 3341 11645 3375 11679
rect 4813 11645 4847 11679
rect 7021 11645 7055 11679
rect 7230 11645 7264 11679
rect 8861 11645 8895 11679
rect 9045 11645 9079 11679
rect 9321 11645 9355 11679
rect 6469 11577 6503 11611
rect 1961 11509 1995 11543
rect 5825 11509 5859 11543
rect 7481 11509 7515 11543
rect 7665 11509 7699 11543
rect 3801 11305 3835 11339
rect 9505 11305 9539 11339
rect 2513 11237 2547 11271
rect 5273 11169 5307 11203
rect 5549 11169 5583 11203
rect 7021 11169 7055 11203
rect 9045 11169 9079 11203
rect 2237 11101 2271 11135
rect 2513 11101 2547 11135
rect 3985 11101 4019 11135
rect 4261 11101 4295 11135
rect 7205 11101 7239 11135
rect 7481 11101 7515 11135
rect 9137 11101 9171 11135
rect 11437 11101 11471 11135
rect 4169 11033 4203 11067
rect 7113 11033 7147 11067
rect 11713 11033 11747 11067
rect 13461 11033 13495 11067
rect 5733 10761 5767 10795
rect 12173 10761 12207 10795
rect 6101 10693 6135 10727
rect 12449 10693 12483 10727
rect 5917 10625 5951 10659
rect 6193 10625 6227 10659
rect 7021 10625 7055 10659
rect 7573 10625 7607 10659
rect 9137 10625 9171 10659
rect 9321 10625 9355 10659
rect 11161 10625 11195 10659
rect 11713 10625 11747 10659
rect 12357 10625 12391 10659
rect 12541 10625 12575 10659
rect 12725 10625 12759 10659
rect 6929 10557 6963 10591
rect 11805 10557 11839 10591
rect 7665 10489 7699 10523
rect 12081 10489 12115 10523
rect 9321 10421 9355 10455
rect 11345 10421 11379 10455
rect 8953 10217 8987 10251
rect 1593 10081 1627 10115
rect 8309 10013 8343 10047
rect 8585 10013 8619 10047
rect 9229 10013 9263 10047
rect 9781 10013 9815 10047
rect 11437 10013 11471 10047
rect 1869 9945 1903 9979
rect 3617 9945 3651 9979
rect 9505 9945 9539 9979
rect 11713 9945 11747 9979
rect 13461 9945 13495 9979
rect 8401 9877 8435 9911
rect 8769 9877 8803 9911
rect 9137 9877 9171 9911
rect 9321 9877 9355 9911
rect 9873 9877 9907 9911
rect 6377 9673 6411 9707
rect 8953 9673 8987 9707
rect 9413 9673 9447 9707
rect 9505 9673 9539 9707
rect 11529 9673 11563 9707
rect 9873 9605 9907 9639
rect 9965 9605 9999 9639
rect 10885 9605 10919 9639
rect 12015 9605 12049 9639
rect 12449 9605 12483 9639
rect 3249 9537 3283 9571
rect 6101 9537 6135 9571
rect 6193 9537 6227 9571
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 7021 9537 7055 9571
rect 8217 9537 8251 9571
rect 9045 9537 9079 9571
rect 10333 9537 10367 9571
rect 10425 9537 10459 9571
rect 10609 9537 10643 9571
rect 10701 9537 10735 9571
rect 11713 9537 11747 9571
rect 11805 9537 11839 9571
rect 11897 9537 11931 9571
rect 12633 9537 12667 9571
rect 12725 9537 12759 9571
rect 12909 9537 12943 9571
rect 13185 9537 13219 9571
rect 1409 9469 1443 9503
rect 1685 9469 1719 9503
rect 3525 9469 3559 9503
rect 5733 9469 5767 9503
rect 5917 9469 5951 9503
rect 8309 9469 8343 9503
rect 8769 9469 8803 9503
rect 10057 9469 10091 9503
rect 12173 9469 12207 9503
rect 8585 9401 8619 9435
rect 12817 9401 12851 9435
rect 13369 9401 13403 9435
rect 3157 9333 3191 9367
rect 4997 9333 5031 9367
rect 12265 9333 12299 9367
rect 2053 9129 2087 9163
rect 3801 9129 3835 9163
rect 5503 9129 5537 9163
rect 6285 9129 6319 9163
rect 6469 9129 6503 9163
rect 7021 9129 7055 9163
rect 8769 9129 8803 9163
rect 9597 9129 9631 9163
rect 1593 9061 1627 9095
rect 4905 9061 4939 9095
rect 5917 9061 5951 9095
rect 7205 9061 7239 9095
rect 2697 8993 2731 9027
rect 4353 8993 4387 9027
rect 5641 8993 5675 9027
rect 7113 8993 7147 9027
rect 9413 8993 9447 9027
rect 9689 8993 9723 9027
rect 1409 8925 1443 8959
rect 1777 8925 1811 8959
rect 1961 8925 1995 8959
rect 3433 8925 3467 8959
rect 4169 8925 4203 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 5365 8925 5399 8959
rect 5825 8925 5859 8959
rect 6561 8925 6595 8959
rect 6837 8925 6871 8959
rect 7297 8925 7331 8959
rect 7389 8925 7423 8959
rect 7941 8925 7975 8959
rect 8033 8925 8067 8959
rect 9045 8925 9079 8959
rect 9321 8925 9355 8959
rect 9873 8925 9907 8959
rect 10149 8925 10183 8959
rect 10333 8925 10367 8959
rect 12265 8925 12299 8959
rect 12541 8925 12575 8959
rect 12633 8925 12667 8959
rect 13185 8925 13219 8959
rect 2513 8857 2547 8891
rect 5733 8857 5767 8891
rect 8217 8857 8251 8891
rect 8401 8857 8435 8891
rect 8953 8857 8987 8891
rect 12725 8857 12759 8891
rect 1869 8789 1903 8823
rect 2421 8789 2455 8823
rect 2973 8789 3007 8823
rect 4261 8789 4295 8823
rect 5181 8789 5215 8823
rect 6285 8789 6319 8823
rect 6653 8789 6687 8823
rect 8493 8789 8527 8823
rect 8585 8789 8619 8823
rect 12081 8789 12115 8823
rect 12449 8789 12483 8823
rect 13369 8789 13403 8823
rect 2513 8585 2547 8619
rect 2973 8585 3007 8619
rect 6193 8585 6227 8619
rect 6653 8585 6687 8619
rect 9045 8585 9079 8619
rect 9137 8585 9171 8619
rect 11345 8585 11379 8619
rect 2237 8517 2271 8551
rect 3893 8517 3927 8551
rect 6377 8517 6411 8551
rect 10977 8517 11011 8551
rect 11193 8517 11227 8551
rect 1409 8449 1443 8483
rect 2881 8449 2915 8483
rect 3709 8449 3743 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 6653 8449 6687 8483
rect 8309 8449 8343 8483
rect 8769 8449 8803 8483
rect 9145 8449 9179 8483
rect 9321 8449 9355 8483
rect 3065 8381 3099 8415
rect 3341 8381 3375 8415
rect 5917 8381 5951 8415
rect 8401 8381 8435 8415
rect 9045 8381 9079 8415
rect 11529 8381 11563 8415
rect 11805 8381 11839 8415
rect 4077 8245 4111 8279
rect 6009 8245 6043 8279
rect 8677 8245 8711 8279
rect 8861 8245 8895 8279
rect 11161 8245 11195 8279
rect 13277 8245 13311 8279
rect 4445 8041 4479 8075
rect 5089 8041 5123 8075
rect 5917 8041 5951 8075
rect 11161 8041 11195 8075
rect 12265 8041 12299 8075
rect 13369 8041 13403 8075
rect 5457 7973 5491 8007
rect 11437 7973 11471 8007
rect 3801 7905 3835 7939
rect 4261 7905 4295 7939
rect 5089 7905 5123 7939
rect 5825 7905 5859 7939
rect 6285 7905 6319 7939
rect 6653 7905 6687 7939
rect 11161 7905 11195 7939
rect 2053 7837 2087 7871
rect 2145 7837 2179 7871
rect 2329 7837 2363 7871
rect 2513 7837 2547 7871
rect 2789 7837 2823 7871
rect 4169 7837 4203 7871
rect 4813 7837 4847 7871
rect 5273 7837 5307 7871
rect 5549 7837 5583 7871
rect 5733 7837 5767 7871
rect 6009 7837 6043 7871
rect 6745 7837 6779 7871
rect 9229 7837 9263 7871
rect 9413 7837 9447 7871
rect 11253 7837 11287 7871
rect 11529 7837 11563 7871
rect 11621 7837 11655 7871
rect 11897 7837 11931 7871
rect 11989 7837 12023 7871
rect 12081 7837 12115 7871
rect 12541 7837 12575 7871
rect 12817 7837 12851 7871
rect 13185 7837 13219 7871
rect 2421 7769 2455 7803
rect 4629 7769 4663 7803
rect 4997 7769 5031 7803
rect 11779 7769 11813 7803
rect 12725 7769 12759 7803
rect 1593 7701 1627 7735
rect 2697 7701 2731 7735
rect 3341 7701 3375 7735
rect 6377 7701 6411 7735
rect 9413 7701 9447 7735
rect 10885 7701 10919 7735
rect 12357 7701 12391 7735
rect 13001 7701 13035 7735
rect 1685 7497 1719 7531
rect 6193 7497 6227 7531
rect 6561 7497 6595 7531
rect 6929 7497 6963 7531
rect 9229 7497 9263 7531
rect 9965 7497 9999 7531
rect 13369 7497 13403 7531
rect 2973 7429 3007 7463
rect 3525 7429 3559 7463
rect 4353 7429 4387 7463
rect 6377 7429 6411 7463
rect 9045 7429 9079 7463
rect 9505 7429 9539 7463
rect 1685 7361 1719 7395
rect 1869 7361 1903 7395
rect 2421 7361 2455 7395
rect 2605 7361 2639 7395
rect 3157 7361 3191 7395
rect 3617 7361 3651 7395
rect 3764 7361 3798 7395
rect 5181 7361 5215 7395
rect 5825 7361 5859 7395
rect 6653 7361 6687 7395
rect 6745 7361 6779 7395
rect 8953 7361 8987 7395
rect 9137 7361 9171 7395
rect 9321 7361 9355 7395
rect 9413 7361 9447 7395
rect 9781 7361 9815 7395
rect 10057 7361 10091 7395
rect 10241 7361 10275 7395
rect 3985 7293 4019 7327
rect 5273 7293 5307 7327
rect 5549 7293 5583 7327
rect 5733 7293 5767 7327
rect 9689 7293 9723 7327
rect 10149 7293 10183 7327
rect 11621 7293 11655 7327
rect 11897 7293 11931 7327
rect 3893 7157 3927 7191
rect 9505 7157 9539 7191
rect 4445 6953 4479 6987
rect 11805 6953 11839 6987
rect 9597 6885 9631 6919
rect 2053 6817 2087 6851
rect 2973 6817 3007 6851
rect 3065 6817 3099 6851
rect 8493 6817 8527 6851
rect 8769 6817 8803 6851
rect 8953 6817 8987 6851
rect 10057 6817 10091 6851
rect 12449 6817 12483 6851
rect 1409 6749 1443 6783
rect 3341 6749 3375 6783
rect 3525 6749 3559 6783
rect 3801 6749 3835 6783
rect 3894 6749 3928 6783
rect 4266 6749 4300 6783
rect 8401 6749 8435 6783
rect 9229 6749 9263 6783
rect 9689 6749 9723 6783
rect 10149 6749 10183 6783
rect 10425 6749 10459 6783
rect 10609 6749 10643 6783
rect 11989 6749 12023 6783
rect 12541 6749 12575 6783
rect 12725 6749 12759 6783
rect 3433 6681 3467 6715
rect 4077 6681 4111 6715
rect 4169 6681 4203 6715
rect 9321 6681 9355 6715
rect 12081 6681 12115 6715
rect 12173 6681 12207 6715
rect 12291 6681 12325 6715
rect 2513 6613 2547 6647
rect 2881 6613 2915 6647
rect 9413 6613 9447 6647
rect 9781 6613 9815 6647
rect 10425 6613 10459 6647
rect 12633 6613 12667 6647
rect 1593 6409 1627 6443
rect 4261 6409 4295 6443
rect 5181 6409 5215 6443
rect 8953 6409 8987 6443
rect 9321 6409 9355 6443
rect 10609 6409 10643 6443
rect 1685 6341 1719 6375
rect 2421 6341 2455 6375
rect 2789 6341 2823 6375
rect 4445 6341 4479 6375
rect 7573 6341 7607 6375
rect 7789 6341 7823 6375
rect 8769 6341 8803 6375
rect 9137 6341 9171 6375
rect 11069 6341 11103 6375
rect 1409 6273 1443 6307
rect 4813 6273 4847 6307
rect 4997 6273 5031 6307
rect 5365 6273 5399 6307
rect 5641 6273 5675 6307
rect 6469 6273 6503 6307
rect 6653 6273 6687 6307
rect 6745 6273 6779 6307
rect 6837 6273 6871 6307
rect 7113 6273 7147 6307
rect 8217 6273 8251 6307
rect 8309 6273 8343 6307
rect 8401 6273 8435 6307
rect 9045 6273 9079 6307
rect 9781 6273 9815 6307
rect 10793 6273 10827 6307
rect 12173 6273 12207 6307
rect 2053 6205 2087 6239
rect 2513 6205 2547 6239
rect 5549 6205 5583 6239
rect 6377 6205 6411 6239
rect 8585 6205 8619 6239
rect 9413 6205 9447 6239
rect 9689 6205 9723 6239
rect 10885 6205 10919 6239
rect 8033 6137 8067 6171
rect 2145 6069 2179 6103
rect 2283 6069 2317 6103
rect 5549 6069 5583 6103
rect 7757 6069 7791 6103
rect 7941 6069 7975 6103
rect 10793 6069 10827 6103
rect 12081 6069 12115 6103
rect 3249 5865 3283 5899
rect 3433 5865 3467 5899
rect 6377 5865 6411 5899
rect 8033 5865 8067 5899
rect 9321 5865 9355 5899
rect 10609 5865 10643 5899
rect 2237 5797 2271 5831
rect 6193 5797 6227 5831
rect 8769 5797 8803 5831
rect 9505 5797 9539 5831
rect 1961 5729 1995 5763
rect 2973 5729 3007 5763
rect 5917 5729 5951 5763
rect 8309 5729 8343 5763
rect 11437 5729 11471 5763
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 2881 5661 2915 5695
rect 3341 5661 3375 5695
rect 3525 5661 3559 5695
rect 5825 5661 5859 5695
rect 6285 5661 6319 5695
rect 6469 5661 6503 5695
rect 6561 5661 6595 5695
rect 6745 5661 6779 5695
rect 7941 5661 7975 5695
rect 8125 5661 8159 5695
rect 8401 5661 8435 5695
rect 9137 5661 9171 5695
rect 9413 5661 9447 5695
rect 9597 5661 9631 5695
rect 10333 5661 10367 5695
rect 10425 5661 10459 5695
rect 10701 5661 10735 5695
rect 11069 5661 11103 5695
rect 11161 5661 11195 5695
rect 8953 5593 8987 5627
rect 10057 5593 10091 5627
rect 10839 5593 10873 5627
rect 10977 5593 11011 5627
rect 11345 5593 11379 5627
rect 11713 5593 11747 5627
rect 13461 5593 13495 5627
rect 1593 5525 1627 5559
rect 6653 5525 6687 5559
rect 10241 5525 10275 5559
rect 1593 5321 1627 5355
rect 2145 5321 2179 5355
rect 3065 5321 3099 5355
rect 5549 5321 5583 5355
rect 7021 5321 7055 5355
rect 11529 5321 11563 5355
rect 12817 5321 12851 5355
rect 2973 5253 3007 5287
rect 12909 5253 12943 5287
rect 1409 5185 1443 5219
rect 4813 5185 4847 5219
rect 4905 5185 4939 5219
rect 5181 5185 5215 5219
rect 5825 5185 5859 5219
rect 6377 5185 6411 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 11897 5185 11931 5219
rect 11989 5185 12023 5219
rect 13185 5185 13219 5219
rect 2237 5117 2271 5151
rect 2421 5117 2455 5151
rect 3157 5117 3191 5151
rect 5089 5117 5123 5151
rect 5273 5117 5307 5151
rect 5917 5117 5951 5151
rect 6193 5117 6227 5151
rect 11713 5117 11747 5151
rect 11805 5117 11839 5151
rect 1777 4981 1811 5015
rect 2605 4981 2639 5015
rect 4997 4981 5031 5015
rect 5181 4981 5215 5015
rect 13369 4981 13403 5015
rect 5825 4777 5859 4811
rect 6101 4777 6135 4811
rect 9505 4777 9539 4811
rect 10609 4777 10643 4811
rect 6745 4709 6779 4743
rect 2973 4641 3007 4675
rect 3157 4641 3191 4675
rect 9229 4641 9263 4675
rect 1501 4573 1535 4607
rect 2053 4573 2087 4607
rect 2881 4573 2915 4607
rect 5733 4573 5767 4607
rect 5917 4573 5951 4607
rect 6561 4573 6595 4607
rect 9137 4573 9171 4607
rect 10241 4573 10275 4607
rect 13461 4573 13495 4607
rect 6285 4505 6319 4539
rect 6469 4505 6503 4539
rect 10425 4505 10459 4539
rect 2513 4437 2547 4471
rect 13277 4437 13311 4471
rect 9045 4233 9079 4267
rect 2605 4165 2639 4199
rect 4353 4165 4387 4199
rect 7113 4165 7147 4199
rect 10149 4165 10183 4199
rect 5825 4097 5859 4131
rect 6561 4097 6595 4131
rect 7021 4097 7055 4131
rect 7297 4097 7331 4131
rect 7665 4097 7699 4131
rect 8585 4097 8619 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10267 4097 10301 4131
rect 2329 4029 2363 4063
rect 5733 4029 5767 4063
rect 6653 4029 6687 4063
rect 6929 4029 6963 4063
rect 7573 4029 7607 4063
rect 9137 4029 9171 4063
rect 9229 4029 9263 4063
rect 10425 4029 10459 4063
rect 6193 3961 6227 3995
rect 8033 3961 8067 3995
rect 7021 3893 7055 3927
rect 8401 3893 8435 3927
rect 8677 3893 8711 3927
rect 9781 3893 9815 3927
rect 1409 3553 1443 3587
rect 1685 3553 1719 3587
rect 5273 3553 5307 3587
rect 7297 3553 7331 3587
rect 9321 3553 9355 3587
rect 9597 3553 9631 3587
rect 11345 3553 11379 3587
rect 3433 3485 3467 3519
rect 7573 3485 7607 3519
rect 7757 3485 7791 3519
rect 7849 3485 7883 3519
rect 5549 3417 5583 3451
rect 7389 3349 7423 3383
rect 6377 3145 6411 3179
rect 7205 3145 7239 3179
rect 10241 3145 10275 3179
rect 10609 3145 10643 3179
rect 2697 3077 2731 3111
rect 6653 3077 6687 3111
rect 7481 3077 7515 3111
rect 8585 3077 8619 3111
rect 10885 3077 10919 3111
rect 2421 3009 2455 3043
rect 6561 3009 6595 3043
rect 6745 3009 6779 3043
rect 6883 3009 6917 3043
rect 7021 3009 7055 3043
rect 10241 3009 10275 3043
rect 10425 3009 10459 3043
rect 4169 2941 4203 2975
rect 8309 2941 8343 2975
rect 10057 2941 10091 2975
rect 7481 2397 7515 2431
rect 8125 2397 8159 2431
rect 8769 2397 8803 2431
rect 7297 2261 7331 2295
rect 7941 2261 7975 2295
rect 8585 2261 8619 2295
<< metal1 >>
rect 1104 14714 13800 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 13800 14714
rect 1104 14640 13800 14662
rect 9674 14560 9680 14612
rect 9732 14600 9738 14612
rect 9861 14603 9919 14609
rect 9861 14600 9873 14603
rect 9732 14572 9873 14600
rect 9732 14560 9738 14572
rect 9861 14569 9873 14572
rect 9907 14569 9919 14603
rect 9861 14563 9919 14569
rect 5810 14424 5816 14476
rect 5868 14464 5874 14476
rect 6733 14467 6791 14473
rect 6733 14464 6745 14467
rect 5868 14436 6745 14464
rect 5868 14424 5874 14436
rect 6733 14433 6745 14436
rect 6779 14433 6791 14467
rect 6733 14427 6791 14433
rect 6181 14399 6239 14405
rect 6181 14365 6193 14399
rect 6227 14396 6239 14399
rect 6362 14396 6368 14408
rect 6227 14368 6368 14396
rect 6227 14365 6239 14368
rect 6181 14359 6239 14365
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 6457 14399 6515 14405
rect 6457 14365 6469 14399
rect 6503 14365 6515 14399
rect 6457 14359 6515 14365
rect 6086 14288 6092 14340
rect 6144 14328 6150 14340
rect 6472 14328 6500 14359
rect 7098 14356 7104 14408
rect 7156 14396 7162 14408
rect 7193 14399 7251 14405
rect 7193 14396 7205 14399
rect 7156 14368 7205 14396
rect 7156 14356 7162 14368
rect 7193 14365 7205 14368
rect 7239 14365 7251 14399
rect 7193 14359 7251 14365
rect 8386 14356 8392 14408
rect 8444 14396 8450 14408
rect 8481 14399 8539 14405
rect 8481 14396 8493 14399
rect 8444 14368 8493 14396
rect 8444 14356 8450 14368
rect 8481 14365 8493 14368
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14396 10103 14399
rect 10318 14396 10324 14408
rect 10091 14368 10324 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 6144 14300 6500 14328
rect 6144 14288 6150 14300
rect 5810 14220 5816 14272
rect 5868 14260 5874 14272
rect 5997 14263 6055 14269
rect 5997 14260 6009 14263
rect 5868 14232 6009 14260
rect 5868 14220 5874 14232
rect 5997 14229 6009 14232
rect 6043 14260 6055 14263
rect 6822 14260 6828 14272
rect 6043 14232 6828 14260
rect 6043 14229 6055 14232
rect 5997 14223 6055 14229
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 7377 14263 7435 14269
rect 7377 14229 7389 14263
rect 7423 14260 7435 14263
rect 7834 14260 7840 14272
rect 7423 14232 7840 14260
rect 7423 14229 7435 14232
rect 7377 14223 7435 14229
rect 7834 14220 7840 14232
rect 7892 14220 7898 14272
rect 8662 14220 8668 14272
rect 8720 14220 8726 14272
rect 1104 14170 13800 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 13800 14170
rect 1104 14096 13800 14118
rect 8018 14056 8024 14068
rect 6380 14028 8024 14056
rect 6380 13929 6408 14028
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 9171 14028 10180 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 6733 13991 6791 13997
rect 6733 13957 6745 13991
rect 6779 13988 6791 13991
rect 7834 13988 7840 14000
rect 6779 13960 7840 13988
rect 6779 13957 6791 13960
rect 6733 13951 6791 13957
rect 7834 13948 7840 13960
rect 7892 13948 7898 14000
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 5442 13812 5448 13864
rect 5500 13812 5506 13864
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 5813 13787 5871 13793
rect 5813 13784 5825 13787
rect 5592 13756 5825 13784
rect 5592 13744 5598 13756
rect 5813 13753 5825 13756
rect 5859 13784 5871 13787
rect 6365 13787 6423 13793
rect 6365 13784 6377 13787
rect 5859 13756 6377 13784
rect 5859 13753 5871 13756
rect 5813 13747 5871 13753
rect 6365 13753 6377 13756
rect 6411 13753 6423 13787
rect 6365 13747 6423 13753
rect 5902 13676 5908 13728
rect 5960 13676 5966 13728
rect 6564 13716 6592 13883
rect 7006 13880 7012 13932
rect 7064 13880 7070 13932
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13920 8999 13923
rect 9140 13920 9168 14019
rect 8987 13892 9168 13920
rect 8987 13889 8999 13892
rect 8941 13883 8999 13889
rect 9398 13880 9404 13932
rect 9456 13920 9462 13932
rect 9493 13923 9551 13929
rect 9493 13920 9505 13923
rect 9456 13892 9505 13920
rect 9456 13880 9462 13892
rect 9493 13889 9505 13892
rect 9539 13889 9551 13923
rect 9493 13883 9551 13889
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13920 9643 13923
rect 9766 13920 9772 13932
rect 9631 13892 9772 13920
rect 9631 13889 9643 13892
rect 9585 13883 9643 13889
rect 9766 13880 9772 13892
rect 9824 13880 9830 13932
rect 10152 13929 10180 14028
rect 10318 14016 10324 14068
rect 10376 14016 10382 14068
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 10686 13920 10692 13932
rect 10183 13892 10692 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 6822 13812 6828 13864
rect 6880 13812 6886 13864
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9677 13815 9735 13821
rect 8478 13744 8484 13796
rect 8536 13784 8542 13796
rect 9692 13784 9720 13815
rect 9950 13812 9956 13864
rect 10008 13812 10014 13864
rect 8536 13756 9720 13784
rect 8536 13744 8542 13756
rect 6733 13719 6791 13725
rect 6733 13716 6745 13719
rect 6564 13688 6745 13716
rect 6733 13685 6745 13688
rect 6779 13716 6791 13719
rect 6914 13716 6920 13728
rect 6779 13688 6920 13716
rect 6779 13685 6791 13688
rect 6733 13679 6791 13685
rect 6914 13676 6920 13688
rect 6972 13676 6978 13728
rect 7190 13676 7196 13728
rect 7248 13676 7254 13728
rect 8754 13676 8760 13728
rect 8812 13716 8818 13728
rect 8849 13719 8907 13725
rect 8849 13716 8861 13719
rect 8812 13688 8861 13716
rect 8812 13676 8818 13688
rect 8849 13685 8861 13688
rect 8895 13685 8907 13719
rect 8849 13679 8907 13685
rect 1104 13626 13800 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 13800 13626
rect 1104 13552 13800 13574
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 5442 13512 5448 13524
rect 5307 13484 5448 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 6254 13515 6312 13521
rect 6254 13512 6266 13515
rect 5960 13484 6266 13512
rect 5960 13472 5966 13484
rect 6254 13481 6266 13484
rect 6300 13481 6312 13515
rect 6254 13475 6312 13481
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7282 13512 7288 13524
rect 7064 13484 7288 13512
rect 7064 13472 7070 13484
rect 7282 13472 7288 13484
rect 7340 13512 7346 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 7340 13484 8953 13512
rect 7340 13472 7346 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 8941 13475 8999 13481
rect 4798 13404 4804 13456
rect 4856 13444 4862 13456
rect 4893 13447 4951 13453
rect 4893 13444 4905 13447
rect 4856 13416 4905 13444
rect 4856 13404 4862 13416
rect 4893 13413 4905 13416
rect 4939 13413 4951 13447
rect 4893 13407 4951 13413
rect 5626 13404 5632 13456
rect 5684 13444 5690 13456
rect 9398 13444 9404 13456
rect 5684 13416 6040 13444
rect 5684 13404 5690 13416
rect 4614 13376 4620 13388
rect 4080 13348 4620 13376
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 4080 13317 4108 13348
rect 4614 13336 4620 13348
rect 4672 13336 4678 13388
rect 4816 13376 4844 13404
rect 5810 13376 5816 13388
rect 4724 13348 4844 13376
rect 5092 13348 5816 13376
rect 4724 13317 4752 13348
rect 5092 13317 5120 13348
rect 5810 13336 5816 13348
rect 5868 13336 5874 13388
rect 6012 13385 6040 13416
rect 7668 13416 9404 13444
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 7668 13376 7696 13416
rect 9398 13404 9404 13416
rect 9456 13404 9462 13456
rect 6043 13348 7696 13376
rect 7745 13379 7803 13385
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 7745 13345 7757 13379
rect 7791 13376 7803 13379
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 7791 13348 8064 13376
rect 7791 13345 7803 13348
rect 7745 13339 7803 13345
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 900 13280 1409 13308
rect 900 13268 906 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 4065 13311 4123 13317
rect 4065 13277 4077 13311
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13277 4583 13311
rect 4525 13271 4583 13277
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 5077 13311 5135 13317
rect 4847 13280 4881 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5077 13277 5089 13311
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 5442 13308 5448 13320
rect 5399 13280 5448 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 4540 13240 4568 13271
rect 4816 13240 4844 13271
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5718 13268 5724 13320
rect 5776 13268 5782 13320
rect 7834 13268 7840 13320
rect 7892 13268 7898 13320
rect 8036 13317 8064 13348
rect 8404 13348 10425 13376
rect 8404 13317 8432 13348
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 10413 13339 10471 13345
rect 10686 13336 10692 13388
rect 10744 13336 10750 13388
rect 8021 13311 8079 13317
rect 8021 13277 8033 13311
rect 8067 13277 8079 13311
rect 8021 13271 8079 13277
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13308 8263 13311
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 8251 13280 8401 13308
rect 8251 13277 8263 13280
rect 8205 13271 8263 13277
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 8662 13308 8668 13320
rect 8619 13280 8668 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 8662 13268 8668 13280
rect 8720 13268 8726 13320
rect 5258 13240 5264 13252
rect 4540 13212 5264 13240
rect 5258 13200 5264 13212
rect 5316 13200 5322 13252
rect 5629 13243 5687 13249
rect 5629 13209 5641 13243
rect 5675 13240 5687 13243
rect 6362 13240 6368 13252
rect 5675 13212 6368 13240
rect 5675 13209 5687 13212
rect 5629 13203 5687 13209
rect 6362 13200 6368 13212
rect 6420 13200 6426 13252
rect 7558 13240 7564 13252
rect 7498 13212 7564 13240
rect 7558 13200 7564 13212
rect 7616 13240 7622 13252
rect 10502 13240 10508 13252
rect 7616 13212 9168 13240
rect 9982 13212 10508 13240
rect 7616 13200 7622 13212
rect 1578 13132 1584 13184
rect 1636 13132 1642 13184
rect 3878 13132 3884 13184
rect 3936 13132 3942 13184
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 5442 13172 5448 13184
rect 4663 13144 5448 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 5902 13132 5908 13184
rect 5960 13132 5966 13184
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 8846 13172 8852 13184
rect 8803 13144 8852 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 8846 13132 8852 13144
rect 8904 13132 8910 13184
rect 9140 13172 9168 13212
rect 10060 13172 10088 13212
rect 10502 13200 10508 13212
rect 10560 13200 10566 13252
rect 9140 13144 10088 13172
rect 1104 13082 13800 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 13800 13082
rect 1104 13008 13800 13030
rect 2682 12968 2688 12980
rect 2608 12940 2688 12968
rect 2608 12909 2636 12940
rect 2682 12928 2688 12940
rect 2740 12968 2746 12980
rect 5626 12968 5632 12980
rect 2740 12940 5632 12968
rect 2740 12928 2746 12940
rect 5626 12928 5632 12940
rect 5684 12928 5690 12980
rect 5997 12971 6055 12977
rect 5997 12937 6009 12971
rect 6043 12968 6055 12971
rect 6086 12968 6092 12980
rect 6043 12940 6092 12968
rect 6043 12937 6055 12940
rect 5997 12931 6055 12937
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 6656 12940 7144 12968
rect 6656 12912 6684 12940
rect 2593 12903 2651 12909
rect 2593 12869 2605 12903
rect 2639 12869 2651 12903
rect 2593 12863 2651 12869
rect 3786 12860 3792 12912
rect 3844 12860 3850 12912
rect 4890 12860 4896 12912
rect 4948 12900 4954 12912
rect 5169 12903 5227 12909
rect 5169 12900 5181 12903
rect 4948 12872 5181 12900
rect 4948 12860 4954 12872
rect 5169 12869 5181 12872
rect 5215 12869 5227 12903
rect 5169 12863 5227 12869
rect 5718 12860 5724 12912
rect 5776 12860 5782 12912
rect 6638 12860 6644 12912
rect 6696 12860 6702 12912
rect 7116 12909 7144 12940
rect 8478 12928 8484 12980
rect 8536 12928 8542 12980
rect 9766 12928 9772 12980
rect 9824 12928 9830 12980
rect 13265 12971 13323 12977
rect 13265 12968 13277 12971
rect 10428 12940 13277 12968
rect 7101 12903 7159 12909
rect 7101 12869 7113 12903
rect 7147 12869 7159 12903
rect 7101 12863 7159 12869
rect 8018 12860 8024 12912
rect 8076 12860 8082 12912
rect 8662 12860 8668 12912
rect 8720 12860 8726 12912
rect 4982 12792 4988 12844
rect 5040 12792 5046 12844
rect 5261 12835 5319 12841
rect 5261 12801 5273 12835
rect 5307 12832 5319 12835
rect 5350 12832 5356 12844
rect 5307 12804 5356 12832
rect 5307 12801 5319 12804
rect 5261 12795 5319 12801
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 5442 12792 5448 12844
rect 5500 12832 5506 12844
rect 5629 12835 5687 12841
rect 5629 12832 5641 12835
rect 5500 12804 5641 12832
rect 5500 12792 5506 12804
rect 5629 12801 5641 12804
rect 5675 12801 5687 12835
rect 5736 12832 5764 12860
rect 5736 12804 6316 12832
rect 5629 12795 5687 12801
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12764 2835 12767
rect 2866 12764 2872 12776
rect 2823 12736 2872 12764
rect 2823 12733 2835 12736
rect 2777 12727 2835 12733
rect 2866 12724 2872 12736
rect 2924 12724 2930 12776
rect 3234 12724 3240 12776
rect 3292 12724 3298 12776
rect 4706 12724 4712 12776
rect 4764 12764 4770 12776
rect 4801 12767 4859 12773
rect 4801 12764 4813 12767
rect 4764 12736 4813 12764
rect 4764 12724 4770 12736
rect 4801 12733 4813 12736
rect 4847 12733 4859 12767
rect 4801 12727 4859 12733
rect 5537 12767 5595 12773
rect 5537 12733 5549 12767
rect 5583 12733 5595 12767
rect 5537 12727 5595 12733
rect 5552 12696 5580 12727
rect 5718 12724 5724 12776
rect 5776 12724 5782 12776
rect 5810 12724 5816 12776
rect 5868 12724 5874 12776
rect 6288 12764 6316 12804
rect 6362 12792 6368 12844
rect 6420 12832 6426 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6420 12804 6837 12832
rect 6420 12792 6426 12804
rect 6825 12801 6837 12804
rect 6871 12832 6883 12835
rect 7006 12832 7012 12844
rect 6871 12804 7012 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 8389 12835 8447 12841
rect 8389 12832 8401 12835
rect 7984 12804 8401 12832
rect 7984 12792 7990 12804
rect 8389 12801 8401 12804
rect 8435 12801 8447 12835
rect 8389 12795 8447 12801
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12832 8631 12835
rect 8680 12832 8708 12860
rect 8619 12804 8708 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8904 12804 8953 12832
rect 8904 12792 8910 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 8941 12795 8999 12801
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12832 10195 12835
rect 10226 12832 10232 12844
rect 10183 12804 10232 12832
rect 10183 12801 10195 12804
rect 10137 12795 10195 12801
rect 10226 12792 10232 12804
rect 10284 12832 10290 12844
rect 10428 12832 10456 12940
rect 13265 12937 13277 12940
rect 13311 12937 13323 12971
rect 13265 12931 13323 12937
rect 10502 12860 10508 12912
rect 10560 12900 10566 12912
rect 10560 12872 12282 12900
rect 10560 12860 10566 12872
rect 10284 12804 10456 12832
rect 10284 12792 10290 12804
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 6288 12736 6561 12764
rect 6549 12733 6561 12736
rect 6595 12764 6607 12767
rect 7561 12767 7619 12773
rect 7561 12764 7573 12767
rect 6595 12736 7573 12764
rect 6595 12733 6607 12736
rect 6549 12727 6607 12733
rect 7561 12733 7573 12736
rect 7607 12733 7619 12767
rect 7561 12727 7619 12733
rect 8662 12724 8668 12776
rect 8720 12724 8726 12776
rect 10042 12724 10048 12776
rect 10100 12724 10106 12776
rect 11517 12767 11575 12773
rect 11517 12764 11529 12767
rect 10152 12736 11529 12764
rect 6454 12696 6460 12708
rect 5552 12668 6460 12696
rect 6454 12656 6460 12668
rect 6512 12656 6518 12708
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 7653 12699 7711 12705
rect 7653 12696 7665 12699
rect 6972 12668 7665 12696
rect 6972 12656 6978 12668
rect 7653 12665 7665 12668
rect 7699 12665 7711 12699
rect 7653 12659 7711 12665
rect 9677 12699 9735 12705
rect 9677 12665 9689 12699
rect 9723 12696 9735 12699
rect 9950 12696 9956 12708
rect 9723 12668 9956 12696
rect 9723 12665 9735 12668
rect 9677 12659 9735 12665
rect 9950 12656 9956 12668
rect 10008 12656 10014 12708
rect 4614 12588 4620 12640
rect 4672 12637 4678 12640
rect 4672 12631 4721 12637
rect 4672 12597 4675 12631
rect 4709 12597 4721 12631
rect 4672 12591 4721 12597
rect 4672 12588 4678 12591
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 7156 12600 7205 12628
rect 7156 12588 7162 12600
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7193 12591 7251 12597
rect 9398 12588 9404 12640
rect 9456 12628 9462 12640
rect 10152 12628 10180 12736
rect 11517 12733 11529 12736
rect 11563 12733 11575 12767
rect 11517 12727 11575 12733
rect 11790 12724 11796 12776
rect 11848 12724 11854 12776
rect 9456 12600 10180 12628
rect 9456 12588 9462 12600
rect 1104 12538 13800 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 13800 12538
rect 1104 12464 13800 12486
rect 3694 12424 3700 12436
rect 2884 12396 3700 12424
rect 2884 12356 2912 12396
rect 3694 12384 3700 12396
rect 3752 12384 3758 12436
rect 4890 12384 4896 12436
rect 4948 12424 4954 12436
rect 5350 12424 5356 12436
rect 4948 12396 5356 12424
rect 4948 12384 4954 12396
rect 5350 12384 5356 12396
rect 5408 12424 5414 12436
rect 5408 12396 6960 12424
rect 5408 12384 5414 12396
rect 2792 12328 2912 12356
rect 3513 12359 3571 12365
rect 1394 12248 1400 12300
rect 1452 12288 1458 12300
rect 2682 12288 2688 12300
rect 1452 12260 2688 12288
rect 1452 12248 1458 12260
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 1762 12180 1768 12232
rect 1820 12180 1826 12232
rect 2792 12138 2820 12328
rect 3513 12325 3525 12359
rect 3559 12356 3571 12359
rect 4154 12356 4160 12368
rect 3559 12328 4160 12356
rect 3559 12325 3571 12328
rect 3513 12319 3571 12325
rect 4154 12316 4160 12328
rect 4212 12356 4218 12368
rect 4982 12356 4988 12368
rect 4212 12328 4988 12356
rect 4212 12316 4218 12328
rect 4982 12316 4988 12328
rect 5040 12316 5046 12368
rect 6932 12356 6960 12396
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 7064 12396 7113 12424
rect 7064 12384 7070 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 7101 12387 7159 12393
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 10042 12424 10048 12436
rect 9447 12396 10048 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 6932 12328 7236 12356
rect 2866 12248 2872 12300
rect 2924 12288 2930 12300
rect 3970 12288 3976 12300
rect 2924 12260 3976 12288
rect 2924 12248 2930 12260
rect 3970 12248 3976 12260
rect 4028 12288 4034 12300
rect 4028 12260 4200 12288
rect 4028 12248 4034 12260
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12220 3387 12223
rect 3375 12192 3464 12220
rect 3375 12189 3387 12192
rect 3329 12183 3387 12189
rect 2958 12112 2964 12164
rect 3016 12152 3022 12164
rect 3436 12152 3464 12192
rect 3510 12180 3516 12232
rect 3568 12220 3574 12232
rect 3881 12223 3939 12229
rect 3881 12220 3893 12223
rect 3568 12192 3893 12220
rect 3568 12180 3574 12192
rect 3881 12189 3893 12192
rect 3927 12189 3939 12223
rect 3881 12183 3939 12189
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 4172 12220 4200 12260
rect 4798 12248 4804 12300
rect 4856 12248 4862 12300
rect 5537 12291 5595 12297
rect 5537 12257 5549 12291
rect 5583 12288 5595 12291
rect 5902 12288 5908 12300
rect 5583 12260 5908 12288
rect 5583 12257 5595 12260
rect 5537 12251 5595 12257
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 6914 12248 6920 12300
rect 6972 12288 6978 12300
rect 7009 12291 7067 12297
rect 7009 12288 7021 12291
rect 6972 12260 7021 12288
rect 6972 12248 6978 12260
rect 7009 12257 7021 12260
rect 7055 12257 7067 12291
rect 7208 12288 7236 12328
rect 7282 12316 7288 12368
rect 7340 12316 7346 12368
rect 10597 12359 10655 12365
rect 10597 12325 10609 12359
rect 10643 12356 10655 12359
rect 11790 12356 11796 12368
rect 10643 12328 11796 12356
rect 10643 12325 10655 12328
rect 10597 12319 10655 12325
rect 11790 12316 11796 12328
rect 11848 12316 11854 12368
rect 9582 12288 9588 12300
rect 7208 12260 9588 12288
rect 7009 12251 7067 12257
rect 5261 12223 5319 12229
rect 5261 12220 5273 12223
rect 4172 12192 5273 12220
rect 5261 12189 5273 12192
rect 5307 12189 5319 12223
rect 7024 12220 7052 12251
rect 7653 12223 7711 12229
rect 7653 12220 7665 12223
rect 7024 12192 7665 12220
rect 5261 12183 5319 12189
rect 7653 12189 7665 12192
rect 7699 12189 7711 12223
rect 7653 12183 7711 12189
rect 7807 12223 7865 12229
rect 7807 12189 7819 12223
rect 7853 12220 7865 12223
rect 8018 12220 8024 12232
rect 7853 12192 8024 12220
rect 7853 12189 7865 12192
rect 7807 12183 7865 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 9324 12229 9352 12260
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 10321 12291 10379 12297
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10870 12288 10876 12300
rect 10367 12260 10876 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 9309 12223 9367 12229
rect 9309 12189 9321 12223
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9490 12180 9496 12232
rect 9548 12180 9554 12232
rect 10226 12180 10232 12232
rect 10284 12180 10290 12232
rect 3016 12124 3464 12152
rect 3016 12112 3022 12124
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 3191 12087 3249 12093
rect 3191 12084 3203 12087
rect 2648 12056 3203 12084
rect 2648 12044 2654 12056
rect 3191 12053 3203 12056
rect 3237 12053 3249 12087
rect 3436 12084 3464 12124
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 4798 12152 4804 12164
rect 3752 12124 4804 12152
rect 3752 12112 3758 12124
rect 4798 12112 4804 12124
rect 4856 12112 4862 12164
rect 5994 12112 6000 12164
rect 6052 12112 6058 12164
rect 7558 12112 7564 12164
rect 7616 12152 7622 12164
rect 7926 12152 7932 12164
rect 7616 12124 7932 12152
rect 7616 12112 7622 12124
rect 7926 12112 7932 12124
rect 7984 12112 7990 12164
rect 6546 12084 6552 12096
rect 3436 12056 6552 12084
rect 3191 12047 3249 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7156 12056 8033 12084
rect 7156 12044 7162 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 1104 11994 13800 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 13800 11994
rect 1104 11920 13800 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1489 11883 1547 11889
rect 1489 11880 1501 11883
rect 1452 11852 1501 11880
rect 1452 11840 1458 11852
rect 1489 11849 1501 11852
rect 1535 11849 1547 11883
rect 1489 11843 1547 11849
rect 1762 11840 1768 11892
rect 1820 11880 1826 11892
rect 2133 11883 2191 11889
rect 2133 11880 2145 11883
rect 1820 11852 2145 11880
rect 1820 11840 1826 11852
rect 2133 11849 2145 11852
rect 2179 11849 2191 11883
rect 2133 11843 2191 11849
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 6914 11880 6920 11892
rect 2648 11852 6920 11880
rect 2648 11840 2654 11852
rect 6914 11840 6920 11852
rect 6972 11840 6978 11892
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7190 11880 7196 11892
rect 7147 11852 7196 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7377 11883 7435 11889
rect 7377 11849 7389 11883
rect 7423 11880 7435 11883
rect 9214 11880 9220 11892
rect 7423 11852 9220 11880
rect 7423 11849 7435 11852
rect 7377 11843 7435 11849
rect 9214 11840 9220 11852
rect 9272 11840 9278 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 10781 11883 10839 11889
rect 10781 11880 10793 11883
rect 9548 11852 10793 11880
rect 9548 11840 9554 11852
rect 10781 11849 10793 11852
rect 10827 11849 10839 11883
rect 10781 11843 10839 11849
rect 1578 11772 1584 11824
rect 1636 11812 1642 11824
rect 1636 11784 2452 11812
rect 1636 11772 1642 11784
rect 1688 11753 1716 11784
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 1765 11747 1823 11753
rect 1765 11713 1777 11747
rect 1811 11713 1823 11747
rect 1765 11707 1823 11713
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 1780 11676 1808 11707
rect 992 11648 1808 11676
rect 992 11636 998 11648
rect 1946 11500 1952 11552
rect 2004 11500 2010 11552
rect 2424 11540 2452 11784
rect 2682 11772 2688 11824
rect 2740 11772 2746 11824
rect 4798 11812 4804 11824
rect 4554 11784 4804 11812
rect 4798 11772 4804 11784
rect 4856 11812 4862 11824
rect 7466 11812 7472 11824
rect 4856 11784 7472 11812
rect 4856 11772 4862 11784
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 9398 11812 9404 11824
rect 8772 11784 9404 11812
rect 2498 11704 2504 11756
rect 2556 11704 2562 11756
rect 2700 11744 2728 11772
rect 3053 11747 3111 11753
rect 3053 11744 3065 11747
rect 2700 11716 3065 11744
rect 3053 11713 3065 11716
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 4890 11704 4896 11756
rect 4948 11744 4954 11756
rect 5442 11744 5448 11756
rect 4948 11716 5448 11744
rect 4948 11704 4954 11716
rect 5442 11704 5448 11716
rect 5500 11744 5506 11756
rect 5500 11716 5672 11744
rect 5500 11704 5506 11716
rect 2777 11679 2835 11685
rect 2777 11645 2789 11679
rect 2823 11676 2835 11679
rect 2958 11676 2964 11688
rect 2823 11648 2964 11676
rect 2823 11645 2835 11648
rect 2777 11639 2835 11645
rect 2958 11636 2964 11648
rect 3016 11636 3022 11688
rect 3329 11679 3387 11685
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 4706 11676 4712 11688
rect 3375 11648 4712 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11676 4859 11679
rect 5350 11676 5356 11688
rect 4847 11648 5356 11676
rect 4847 11645 4859 11648
rect 4801 11639 4859 11645
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5644 11676 5672 11716
rect 5718 11704 5724 11756
rect 5776 11704 5782 11756
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11744 5963 11747
rect 6365 11747 6423 11753
rect 6365 11744 6377 11747
rect 5951 11716 6377 11744
rect 5951 11713 5963 11716
rect 5905 11707 5963 11713
rect 6365 11713 6377 11716
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 6733 11747 6791 11753
rect 6733 11713 6745 11747
rect 6779 11744 6791 11747
rect 6914 11744 6920 11756
rect 6779 11716 6920 11744
rect 6779 11713 6791 11716
rect 6733 11707 6791 11713
rect 5920 11676 5948 11707
rect 5644 11648 5948 11676
rect 6380 11676 6408 11707
rect 6914 11704 6920 11716
rect 6972 11744 6978 11756
rect 7558 11744 7564 11756
rect 6972 11716 7564 11744
rect 6972 11704 6978 11716
rect 7558 11704 7564 11716
rect 7616 11744 7622 11756
rect 7653 11747 7711 11753
rect 7653 11744 7665 11747
rect 7616 11716 7665 11744
rect 7616 11704 7622 11716
rect 7653 11713 7665 11716
rect 7699 11713 7711 11747
rect 7653 11707 7711 11713
rect 7834 11704 7840 11756
rect 7892 11704 7898 11756
rect 8772 11753 8800 11784
rect 9398 11772 9404 11784
rect 9456 11772 9462 11824
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11713 8815 11747
rect 8757 11707 8815 11713
rect 10410 11704 10416 11756
rect 10468 11704 10474 11756
rect 7006 11676 7012 11688
rect 6380 11648 7012 11676
rect 7006 11636 7012 11648
rect 7064 11636 7070 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7218 11679 7276 11685
rect 7218 11676 7230 11679
rect 7156 11648 7230 11676
rect 7156 11636 7162 11648
rect 7218 11645 7230 11648
rect 7264 11645 7276 11679
rect 7218 11639 7276 11645
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11676 8907 11679
rect 9033 11679 9091 11685
rect 9033 11676 9045 11679
rect 8895 11648 9045 11676
rect 8895 11645 8907 11648
rect 8849 11639 8907 11645
rect 9033 11645 9045 11648
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9306 11636 9312 11688
rect 9364 11636 9370 11688
rect 6454 11568 6460 11620
rect 6512 11608 6518 11620
rect 6512 11580 7696 11608
rect 6512 11568 6518 11580
rect 4706 11540 4712 11552
rect 2424 11512 4712 11540
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 5534 11500 5540 11552
rect 5592 11540 5598 11552
rect 5813 11543 5871 11549
rect 5813 11540 5825 11543
rect 5592 11512 5825 11540
rect 5592 11500 5598 11512
rect 5813 11509 5825 11512
rect 5859 11509 5871 11543
rect 5813 11503 5871 11509
rect 7469 11543 7527 11549
rect 7469 11509 7481 11543
rect 7515 11540 7527 11543
rect 7558 11540 7564 11552
rect 7515 11512 7564 11540
rect 7515 11509 7527 11512
rect 7469 11503 7527 11509
rect 7558 11500 7564 11512
rect 7616 11500 7622 11552
rect 7668 11549 7696 11580
rect 7653 11543 7711 11549
rect 7653 11509 7665 11543
rect 7699 11509 7711 11543
rect 7653 11503 7711 11509
rect 1104 11450 13800 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 13800 11450
rect 1104 11376 13800 11398
rect 3234 11296 3240 11348
rect 3292 11336 3298 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3292 11308 3801 11336
rect 3292 11296 3298 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 4764 11308 6592 11336
rect 4764 11296 4770 11308
rect 2501 11271 2559 11277
rect 2501 11237 2513 11271
rect 2547 11268 2559 11271
rect 3510 11268 3516 11280
rect 2547 11240 3516 11268
rect 2547 11237 2559 11240
rect 2501 11231 2559 11237
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 3970 11228 3976 11280
rect 4028 11228 4034 11280
rect 6564 11268 6592 11308
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9493 11339 9551 11345
rect 9493 11336 9505 11339
rect 9364 11308 9505 11336
rect 9364 11296 9370 11308
rect 9493 11305 9505 11308
rect 9539 11305 9551 11339
rect 9493 11299 9551 11305
rect 11146 11268 11152 11280
rect 6564 11240 11152 11268
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 3234 11160 3240 11212
rect 3292 11200 3298 11212
rect 3988 11200 4016 11228
rect 5261 11203 5319 11209
rect 5261 11200 5273 11203
rect 3292 11172 5273 11200
rect 3292 11160 3298 11172
rect 5261 11169 5273 11172
rect 5307 11169 5319 11203
rect 5261 11163 5319 11169
rect 5534 11160 5540 11212
rect 5592 11160 5598 11212
rect 7009 11203 7067 11209
rect 7009 11169 7021 11203
rect 7055 11200 7067 11203
rect 7055 11172 7512 11200
rect 7055 11169 7067 11172
rect 7009 11163 7067 11169
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 2004 11104 2237 11132
rect 2004 11092 2010 11104
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2498 11092 2504 11144
rect 2556 11092 2562 11144
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4062 11132 4068 11144
rect 4019 11104 4068 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11132 4307 11135
rect 4706 11132 4712 11144
rect 4295 11104 4712 11132
rect 4295 11101 4307 11104
rect 4249 11095 4307 11101
rect 4706 11092 4712 11104
rect 4764 11092 4770 11144
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 7484 11141 7512 11172
rect 9030 11160 9036 11212
rect 9088 11160 9094 11212
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11132 7527 11135
rect 8018 11132 8024 11144
rect 7515 11104 8024 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9490 11132 9496 11144
rect 9171 11104 9496 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9490 11092 9496 11104
rect 9548 11092 9554 11144
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 4614 11064 4620 11076
rect 4203 11036 4620 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 4614 11024 4620 11036
rect 4672 11024 4678 11076
rect 5534 11024 5540 11076
rect 5592 11064 5598 11076
rect 5994 11064 6000 11076
rect 5592 11036 6000 11064
rect 5592 11024 5598 11036
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 7101 11067 7159 11073
rect 7101 11033 7113 11067
rect 7147 11064 7159 11067
rect 7834 11064 7840 11076
rect 7147 11036 7840 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 7834 11024 7840 11036
rect 7892 11064 7898 11076
rect 7892 11036 11100 11064
rect 7892 11024 7898 11036
rect 11072 10996 11100 11036
rect 11698 11024 11704 11076
rect 11756 11024 11762 11076
rect 12710 11024 12716 11076
rect 12768 11024 12774 11076
rect 13170 11024 13176 11076
rect 13228 11064 13234 11076
rect 13449 11067 13507 11073
rect 13449 11064 13461 11067
rect 13228 11036 13461 11064
rect 13228 11024 13234 11036
rect 13449 11033 13461 11036
rect 13495 11033 13507 11067
rect 13449 11027 13507 11033
rect 11882 10996 11888 11008
rect 11072 10968 11888 10996
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 1104 10906 13800 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 13800 10906
rect 1104 10832 13800 10854
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 4614 10792 4620 10804
rect 3936 10764 4620 10792
rect 3936 10752 3942 10764
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 5718 10752 5724 10804
rect 5776 10752 5782 10804
rect 7098 10792 7104 10804
rect 5920 10764 7104 10792
rect 5920 10665 5948 10764
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 11698 10752 11704 10804
rect 11756 10792 11762 10804
rect 12161 10795 12219 10801
rect 12161 10792 12173 10795
rect 11756 10764 12173 10792
rect 11756 10752 11762 10764
rect 12161 10761 12173 10764
rect 12207 10761 12219 10795
rect 12161 10755 12219 10761
rect 6089 10727 6147 10733
rect 6089 10693 6101 10727
rect 6135 10724 6147 10727
rect 6362 10724 6368 10736
rect 6135 10696 6368 10724
rect 6135 10693 6147 10696
rect 6089 10687 6147 10693
rect 6362 10684 6368 10696
rect 6420 10724 6426 10736
rect 12437 10727 12495 10733
rect 12437 10724 12449 10727
rect 6420 10696 7052 10724
rect 6420 10684 6426 10696
rect 7024 10665 7052 10696
rect 11716 10696 12449 10724
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 5905 10619 5963 10625
rect 6181 10659 6239 10665
rect 6181 10625 6193 10659
rect 6227 10656 6239 10659
rect 7009 10659 7067 10665
rect 6227 10628 6960 10656
rect 6227 10625 6239 10628
rect 6181 10619 6239 10625
rect 6932 10600 6960 10628
rect 7009 10625 7021 10659
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7558 10616 7564 10668
rect 7616 10616 7622 10668
rect 9122 10616 9128 10668
rect 9180 10616 9186 10668
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9582 10656 9588 10668
rect 9355 10628 9588 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 11146 10616 11152 10668
rect 11204 10616 11210 10668
rect 11716 10665 11744 10696
rect 12437 10693 12449 10696
rect 12483 10724 12495 10727
rect 13170 10724 13176 10736
rect 12483 10696 13176 10724
rect 12483 10693 12495 10696
rect 12437 10687 12495 10693
rect 13170 10684 13176 10696
rect 13228 10684 13234 10736
rect 11701 10659 11759 10665
rect 11701 10625 11713 10659
rect 11747 10625 11759 10659
rect 11701 10619 11759 10625
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 8570 10548 8576 10600
rect 8628 10588 8634 10600
rect 11716 10588 11744 10619
rect 11882 10616 11888 10668
rect 11940 10656 11946 10668
rect 12250 10656 12256 10668
rect 11940 10628 12256 10656
rect 11940 10616 11946 10628
rect 12250 10616 12256 10628
rect 12308 10656 12314 10668
rect 12345 10659 12403 10665
rect 12345 10656 12357 10659
rect 12308 10628 12357 10656
rect 12308 10616 12314 10628
rect 12345 10625 12357 10628
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10625 12587 10659
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 12529 10619 12587 10625
rect 12636 10628 12725 10656
rect 8628 10560 11744 10588
rect 8628 10548 8634 10560
rect 11790 10548 11796 10600
rect 11848 10548 11854 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12544 10588 12572 10619
rect 12492 10560 12572 10588
rect 12492 10548 12498 10560
rect 7653 10523 7711 10529
rect 7653 10489 7665 10523
rect 7699 10520 7711 10523
rect 11882 10520 11888 10532
rect 7699 10492 11888 10520
rect 7699 10489 7711 10492
rect 7653 10483 7711 10489
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10520 12127 10523
rect 12636 10520 12664 10628
rect 12713 10625 12725 10628
rect 12759 10625 12771 10659
rect 12713 10619 12771 10625
rect 12115 10492 12664 10520
rect 12115 10489 12127 10492
rect 12069 10483 12127 10489
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9950 10452 9956 10464
rect 9355 10424 9956 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 11333 10455 11391 10461
rect 11333 10421 11345 10455
rect 11379 10452 11391 10455
rect 11422 10452 11428 10464
rect 11379 10424 11428 10452
rect 11379 10421 11391 10424
rect 11333 10415 11391 10421
rect 11422 10412 11428 10424
rect 11480 10412 11486 10464
rect 11900 10452 11928 10480
rect 12342 10452 12348 10464
rect 11900 10424 12348 10452
rect 12342 10412 12348 10424
rect 12400 10412 12406 10464
rect 1104 10362 13800 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 13800 10362
rect 1104 10288 13800 10310
rect 8941 10251 8999 10257
rect 8941 10217 8953 10251
rect 8987 10248 8999 10251
rect 9030 10248 9036 10260
rect 8987 10220 9036 10248
rect 8987 10217 8999 10220
rect 8941 10211 8999 10217
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 1394 10072 1400 10124
rect 1452 10112 1458 10124
rect 1581 10115 1639 10121
rect 1581 10112 1593 10115
rect 1452 10084 1593 10112
rect 1452 10072 1458 10084
rect 1581 10081 1593 10084
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 3694 10044 3700 10056
rect 2990 10016 3700 10044
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 8570 10004 8576 10056
rect 8628 10004 8634 10056
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 9769 10047 9827 10053
rect 9769 10044 9781 10047
rect 9272 10016 9781 10044
rect 9272 10004 9278 10016
rect 9769 10013 9781 10016
rect 9815 10013 9827 10047
rect 9769 10007 9827 10013
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 1854 9936 1860 9988
rect 1912 9936 1918 9988
rect 3605 9979 3663 9985
rect 3605 9945 3617 9979
rect 3651 9945 3663 9979
rect 3605 9939 3663 9945
rect 3620 9908 3648 9939
rect 9490 9936 9496 9988
rect 9548 9936 9554 9988
rect 11698 9936 11704 9988
rect 11756 9936 11762 9988
rect 12710 9936 12716 9988
rect 12768 9936 12774 9988
rect 13078 9936 13084 9988
rect 13136 9976 13142 9988
rect 13449 9979 13507 9985
rect 13449 9976 13461 9979
rect 13136 9948 13461 9976
rect 13136 9936 13142 9948
rect 13449 9945 13461 9948
rect 13495 9945 13507 9979
rect 13449 9939 13507 9945
rect 3694 9908 3700 9920
rect 3620 9880 3700 9908
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 8386 9868 8392 9920
rect 8444 9868 8450 9920
rect 8754 9868 8760 9920
rect 8812 9868 8818 9920
rect 9030 9868 9036 9920
rect 9088 9908 9094 9920
rect 9125 9911 9183 9917
rect 9125 9908 9137 9911
rect 9088 9880 9137 9908
rect 9088 9868 9094 9880
rect 9125 9877 9137 9880
rect 9171 9877 9183 9911
rect 9125 9871 9183 9877
rect 9306 9868 9312 9920
rect 9364 9868 9370 9920
rect 9861 9911 9919 9917
rect 9861 9877 9873 9911
rect 9907 9908 9919 9911
rect 10318 9908 10324 9920
rect 9907 9880 10324 9908
rect 9907 9877 9919 9880
rect 9861 9871 9919 9877
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 1104 9818 13800 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 13800 9818
rect 1104 9744 13800 9766
rect 6362 9664 6368 9716
rect 6420 9664 6426 9716
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 8941 9707 8999 9713
rect 8941 9704 8953 9707
rect 8812 9676 8953 9704
rect 8812 9664 8818 9676
rect 8941 9673 8953 9676
rect 8987 9673 8999 9707
rect 8941 9667 8999 9673
rect 9306 9664 9312 9716
rect 9364 9704 9370 9716
rect 9401 9707 9459 9713
rect 9401 9704 9413 9707
rect 9364 9676 9413 9704
rect 9364 9664 9370 9676
rect 9401 9673 9413 9676
rect 9447 9673 9459 9707
rect 9401 9667 9459 9673
rect 9490 9664 9496 9716
rect 9548 9664 9554 9716
rect 11517 9707 11575 9713
rect 11517 9673 11529 9707
rect 11563 9704 11575 9707
rect 11698 9704 11704 9716
rect 11563 9676 11704 9704
rect 11563 9673 11575 9676
rect 11517 9667 11575 9673
rect 11698 9664 11704 9676
rect 11756 9664 11762 9716
rect 12158 9704 12164 9716
rect 11992 9676 12164 9704
rect 3970 9636 3976 9648
rect 2898 9608 3976 9636
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6604 9608 7972 9636
rect 6604 9596 6610 9608
rect 7944 9580 7972 9608
rect 8570 9596 8576 9648
rect 8628 9636 8634 9648
rect 8628 9608 9168 9636
rect 8628 9596 8634 9608
rect 3234 9528 3240 9580
rect 3292 9528 3298 9580
rect 6086 9528 6092 9580
rect 6144 9528 6150 9580
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6270 9568 6276 9580
rect 6227 9540 6276 9568
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6270 9528 6276 9540
rect 6328 9528 6334 9580
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 6641 9571 6699 9577
rect 6641 9568 6653 9571
rect 6512 9540 6653 9568
rect 6512 9528 6518 9540
rect 6641 9537 6653 9540
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 6733 9531 6791 9537
rect 1397 9503 1455 9509
rect 1397 9469 1409 9503
rect 1443 9500 1455 9503
rect 1443 9472 1532 9500
rect 1443 9469 1455 9472
rect 1397 9463 1455 9469
rect 1504 9364 1532 9472
rect 1670 9460 1676 9512
rect 1728 9460 1734 9512
rect 2222 9460 2228 9512
rect 2280 9500 2286 9512
rect 3252 9500 3280 9528
rect 2280 9472 3280 9500
rect 2280 9460 2286 9472
rect 3510 9460 3516 9512
rect 3568 9460 3574 9512
rect 3970 9460 3976 9512
rect 4028 9500 4034 9512
rect 5534 9500 5540 9512
rect 4028 9472 5540 9500
rect 4028 9460 4034 9472
rect 5534 9460 5540 9472
rect 5592 9460 5598 9512
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9500 5779 9503
rect 5810 9500 5816 9512
rect 5767 9472 5816 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 5810 9460 5816 9472
rect 5868 9460 5874 9512
rect 5905 9503 5963 9509
rect 5905 9469 5917 9503
rect 5951 9500 5963 9503
rect 6748 9500 6776 9531
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 7006 9528 7012 9580
rect 7064 9528 7070 9580
rect 7926 9528 7932 9580
rect 7984 9568 7990 9580
rect 8205 9571 8263 9577
rect 8205 9568 8217 9571
rect 7984 9540 8217 9568
rect 7984 9528 7990 9540
rect 8205 9537 8217 9540
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 9140 9568 9168 9608
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9640 9608 9873 9636
rect 9640 9596 9646 9608
rect 9861 9605 9873 9608
rect 9907 9605 9919 9639
rect 9861 9599 9919 9605
rect 9950 9596 9956 9648
rect 10008 9596 10014 9648
rect 10870 9596 10876 9648
rect 10928 9596 10934 9648
rect 11992 9645 12020 9676
rect 12158 9664 12164 9676
rect 12216 9664 12222 9716
rect 11992 9639 12061 9645
rect 11992 9608 12015 9639
rect 12003 9605 12015 9608
rect 12049 9605 12061 9639
rect 12437 9639 12495 9645
rect 12437 9636 12449 9639
rect 12003 9599 12061 9605
rect 12176 9608 12449 9636
rect 9140 9540 10272 9568
rect 9033 9531 9091 9537
rect 5951 9472 6776 9500
rect 5951 9469 5963 9472
rect 5905 9463 5963 9469
rect 8294 9460 8300 9512
rect 8352 9460 8358 9512
rect 8754 9460 8760 9512
rect 8812 9460 8818 9512
rect 9048 9500 9076 9531
rect 9858 9500 9864 9512
rect 9048 9472 9864 9500
rect 8573 9435 8631 9441
rect 8573 9401 8585 9435
rect 8619 9432 8631 9435
rect 9048 9432 9076 9472
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 10042 9460 10048 9512
rect 10100 9460 10106 9512
rect 10244 9500 10272 9540
rect 10318 9528 10324 9580
rect 10376 9528 10382 9580
rect 10413 9571 10471 9577
rect 10413 9537 10425 9571
rect 10459 9537 10471 9571
rect 10413 9531 10471 9537
rect 10428 9500 10456 9531
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 10686 9528 10692 9580
rect 10744 9528 10750 9580
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 10244 9472 10456 9500
rect 8619 9404 9076 9432
rect 8619 9401 8631 9404
rect 8573 9395 8631 9401
rect 2222 9364 2228 9376
rect 1504 9336 2228 9364
rect 2222 9324 2228 9336
rect 2280 9324 2286 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 4798 9364 4804 9376
rect 3191 9336 4804 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 4798 9324 4804 9336
rect 4856 9324 4862 9376
rect 4985 9367 5043 9373
rect 4985 9333 4997 9367
rect 5031 9364 5043 9367
rect 5534 9364 5540 9376
rect 5031 9336 5540 9364
rect 5031 9333 5043 9336
rect 4985 9327 5043 9333
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 8110 9364 8116 9376
rect 5960 9336 8116 9364
rect 5960 9324 5966 9336
rect 8110 9324 8116 9336
rect 8168 9324 8174 9376
rect 11716 9364 11744 9531
rect 11790 9528 11796 9580
rect 11848 9528 11854 9580
rect 11882 9528 11888 9580
rect 11940 9528 11946 9580
rect 11808 9432 11836 9528
rect 12176 9512 12204 9608
rect 12437 9605 12449 9608
rect 12483 9636 12495 9639
rect 13078 9636 13084 9648
rect 12483 9608 13084 9636
rect 12483 9605 12495 9608
rect 12437 9599 12495 9605
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 12912 9577 12940 9608
rect 13078 9596 13084 9608
rect 13136 9596 13142 9648
rect 12713 9571 12771 9577
rect 12713 9568 12725 9571
rect 12676 9540 12725 9568
rect 12676 9528 12682 9540
rect 12713 9537 12725 9540
rect 12759 9537 12771 9571
rect 12713 9531 12771 9537
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9537 12955 9571
rect 12897 9531 12955 9537
rect 13170 9528 13176 9580
rect 13228 9528 13234 9580
rect 12158 9460 12164 9512
rect 12216 9460 12222 9512
rect 12805 9435 12863 9441
rect 12805 9432 12817 9435
rect 11808 9404 12817 9432
rect 12805 9401 12817 9404
rect 12851 9401 12863 9435
rect 12805 9395 12863 9401
rect 13354 9392 13360 9444
rect 13412 9392 13418 9444
rect 12253 9367 12311 9373
rect 12253 9364 12265 9367
rect 11716 9336 12265 9364
rect 12253 9333 12265 9336
rect 12299 9333 12311 9367
rect 12253 9327 12311 9333
rect 1104 9274 13800 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 13800 9274
rect 1104 9200 13800 9222
rect 1854 9120 1860 9172
rect 1912 9160 1918 9172
rect 2041 9163 2099 9169
rect 2041 9160 2053 9163
rect 1912 9132 2053 9160
rect 1912 9120 1918 9132
rect 2041 9129 2053 9132
rect 2087 9129 2099 9163
rect 2041 9123 2099 9129
rect 3510 9120 3516 9172
rect 3568 9160 3574 9172
rect 3789 9163 3847 9169
rect 3789 9160 3801 9163
rect 3568 9132 3801 9160
rect 3568 9120 3574 9132
rect 3789 9129 3801 9132
rect 3835 9129 3847 9163
rect 5491 9163 5549 9169
rect 5491 9160 5503 9163
rect 3789 9123 3847 9129
rect 4908 9132 5503 9160
rect 1581 9095 1639 9101
rect 1581 9061 1593 9095
rect 1627 9092 1639 9095
rect 2314 9092 2320 9104
rect 1627 9064 2320 9092
rect 1627 9061 1639 9064
rect 1581 9055 1639 9061
rect 2314 9052 2320 9064
rect 2372 9092 2378 9104
rect 2372 9064 4200 9092
rect 2372 9052 2378 9064
rect 2590 9024 2596 9036
rect 1964 8996 2596 9024
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 1964 8965 1992 8996
rect 2590 8984 2596 8996
rect 2648 8984 2654 9036
rect 2682 8984 2688 9036
rect 2740 8984 2746 9036
rect 4172 8965 4200 9064
rect 4706 9052 4712 9104
rect 4764 9052 4770 9104
rect 4908 9101 4936 9132
rect 5491 9129 5503 9132
rect 5537 9160 5549 9163
rect 5626 9160 5632 9172
rect 5537 9132 5632 9160
rect 5537 9129 5549 9132
rect 5491 9123 5549 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 6144 9132 6285 9160
rect 6144 9120 6150 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 6273 9123 6331 9129
rect 6454 9120 6460 9172
rect 6512 9120 6518 9172
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7009 9163 7067 9169
rect 7009 9160 7021 9163
rect 6880 9132 7021 9160
rect 6880 9120 6886 9132
rect 7009 9129 7021 9132
rect 7055 9129 7067 9163
rect 7009 9123 7067 9129
rect 8754 9120 8760 9172
rect 8812 9120 8818 9172
rect 9585 9163 9643 9169
rect 9585 9129 9597 9163
rect 9631 9160 9643 9163
rect 10042 9160 10048 9172
rect 9631 9132 10048 9160
rect 9631 9129 9643 9132
rect 9585 9123 9643 9129
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 12158 9160 12164 9172
rect 11296 9132 12164 9160
rect 11296 9120 11302 9132
rect 12158 9120 12164 9132
rect 12216 9120 12222 9172
rect 4893 9095 4951 9101
rect 4893 9061 4905 9095
rect 4939 9061 4951 9095
rect 4893 9055 4951 9061
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 5905 9095 5963 9101
rect 5905 9092 5917 9095
rect 5868 9064 5917 9092
rect 5868 9052 5874 9064
rect 5905 9061 5917 9064
rect 5951 9092 5963 9095
rect 6178 9092 6184 9104
rect 5951 9064 6184 9092
rect 5951 9061 5963 9064
rect 5905 9055 5963 9061
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 7193 9095 7251 9101
rect 7193 9092 7205 9095
rect 6288 9064 7205 9092
rect 4338 8984 4344 9036
rect 4396 9024 4402 9036
rect 4724 9024 4752 9052
rect 6288 9036 6316 9064
rect 7193 9061 7205 9064
rect 7239 9061 7251 9095
rect 8938 9092 8944 9104
rect 7193 9055 7251 9061
rect 7300 9064 8944 9092
rect 4396 8996 4752 9024
rect 5629 9027 5687 9033
rect 4396 8984 4402 8996
rect 5629 8993 5641 9027
rect 5675 9024 5687 9027
rect 5718 9024 5724 9036
rect 5675 8996 5724 9024
rect 5675 8993 5687 8996
rect 5629 8987 5687 8993
rect 5718 8984 5724 8996
rect 5776 9024 5782 9036
rect 5776 8996 6040 9024
rect 5776 8984 5782 8996
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 3421 8959 3479 8965
rect 3421 8956 3433 8959
rect 1949 8919 2007 8925
rect 2424 8928 3433 8956
rect 2424 8832 2452 8928
rect 3421 8925 3433 8928
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4614 8956 4620 8968
rect 4203 8928 4620 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8956 4767 8959
rect 4798 8956 4804 8968
rect 4755 8928 4804 8956
rect 4755 8925 4767 8928
rect 4709 8919 4767 8925
rect 4798 8916 4804 8928
rect 4856 8916 4862 8968
rect 4985 8959 5043 8965
rect 4985 8925 4997 8959
rect 5031 8925 5043 8959
rect 4985 8919 5043 8925
rect 2501 8891 2559 8897
rect 2501 8857 2513 8891
rect 2547 8888 2559 8891
rect 3694 8888 3700 8900
rect 2547 8860 3700 8888
rect 2547 8857 2559 8860
rect 2501 8851 2559 8857
rect 3694 8848 3700 8860
rect 3752 8848 3758 8900
rect 4338 8888 4344 8900
rect 4172 8860 4344 8888
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8820 1915 8823
rect 2130 8820 2136 8832
rect 1903 8792 2136 8820
rect 1903 8789 1915 8792
rect 1857 8783 1915 8789
rect 2130 8780 2136 8792
rect 2188 8780 2194 8832
rect 2406 8780 2412 8832
rect 2464 8780 2470 8832
rect 2958 8780 2964 8832
rect 3016 8780 3022 8832
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 4172 8820 4200 8860
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 5000 8888 5028 8919
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8956 5871 8959
rect 5902 8956 5908 8968
rect 5859 8928 5908 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 6012 8956 6040 8996
rect 6270 8984 6276 9036
rect 6328 8984 6334 9036
rect 6730 9024 6736 9036
rect 6380 8996 6736 9024
rect 6380 8956 6408 8996
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 7101 9027 7159 9033
rect 7101 9024 7113 9027
rect 6932 8996 7113 9024
rect 6012 8928 6408 8956
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 5721 8891 5779 8897
rect 5000 8860 5580 8888
rect 5552 8832 5580 8860
rect 5721 8857 5733 8891
rect 5767 8888 5779 8891
rect 6362 8888 6368 8900
rect 5767 8860 6368 8888
rect 5767 8857 5779 8860
rect 5721 8851 5779 8857
rect 6362 8848 6368 8860
rect 6420 8888 6426 8900
rect 6564 8888 6592 8919
rect 6638 8916 6644 8968
rect 6696 8956 6702 8968
rect 6825 8959 6883 8965
rect 6825 8956 6837 8959
rect 6696 8928 6837 8956
rect 6696 8916 6702 8928
rect 6825 8925 6837 8928
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 6420 8860 6592 8888
rect 6420 8848 6426 8860
rect 6730 8848 6736 8900
rect 6788 8888 6794 8900
rect 6932 8888 6960 8996
rect 7101 8993 7113 8996
rect 7147 9024 7159 9027
rect 7300 9024 7328 9064
rect 8938 9052 8944 9064
rect 8996 9092 9002 9104
rect 8996 9064 10364 9092
rect 8996 9052 9002 9064
rect 7147 8996 7328 9024
rect 7147 8993 7159 8996
rect 7101 8987 7159 8993
rect 8386 8984 8392 9036
rect 8444 8984 8450 9036
rect 8662 8984 8668 9036
rect 8720 9024 8726 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 8720 8996 9413 9024
rect 8720 8984 8726 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 7377 8959 7435 8965
rect 7377 8925 7389 8959
rect 7423 8925 7435 8959
rect 7377 8919 7435 8925
rect 6788 8860 6960 8888
rect 6788 8848 6794 8860
rect 3108 8792 4200 8820
rect 4249 8823 4307 8829
rect 3108 8780 3114 8792
rect 4249 8789 4261 8823
rect 4295 8820 4307 8823
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 4295 8792 5181 8820
rect 4295 8789 4307 8792
rect 4249 8783 4307 8789
rect 5169 8789 5181 8792
rect 5215 8820 5227 8823
rect 5350 8820 5356 8832
rect 5215 8792 5356 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5534 8780 5540 8832
rect 5592 8780 5598 8832
rect 6270 8780 6276 8832
rect 6328 8780 6334 8832
rect 6454 8780 6460 8832
rect 6512 8820 6518 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 6512 8792 6653 8820
rect 6512 8780 6518 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 6641 8783 6699 8789
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 7300 8820 7328 8919
rect 7392 8888 7420 8919
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 8021 8959 8079 8965
rect 8021 8925 8033 8959
rect 8067 8956 8079 8959
rect 8404 8956 8432 8984
rect 8754 8956 8760 8968
rect 8067 8928 8760 8956
rect 8067 8925 8079 8928
rect 8021 8919 8079 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 9033 8959 9091 8965
rect 9033 8956 9045 8959
rect 8904 8928 9045 8956
rect 8904 8916 8910 8928
rect 9033 8925 9045 8928
rect 9079 8925 9091 8959
rect 9033 8919 9091 8925
rect 8202 8888 8208 8900
rect 7392 8860 8208 8888
rect 8202 8848 8208 8860
rect 8260 8848 8266 8900
rect 8389 8891 8447 8897
rect 8389 8857 8401 8891
rect 8435 8888 8447 8891
rect 8938 8888 8944 8900
rect 8435 8860 8944 8888
rect 8435 8857 8447 8860
rect 8389 8851 8447 8857
rect 8938 8848 8944 8860
rect 8996 8848 9002 8900
rect 9048 8888 9076 8919
rect 9122 8916 9128 8968
rect 9180 8956 9186 8968
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 9180 8928 9321 8956
rect 9180 8916 9186 8928
rect 9309 8925 9321 8928
rect 9355 8925 9367 8959
rect 9416 8956 9444 8987
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9677 9027 9735 9033
rect 9677 9024 9689 9027
rect 9640 8996 9689 9024
rect 9640 8984 9646 8996
rect 9677 8993 9689 8996
rect 9723 8993 9735 9027
rect 9677 8987 9735 8993
rect 10336 8965 10364 9064
rect 9861 8959 9919 8965
rect 9861 8956 9873 8959
rect 9416 8928 9873 8956
rect 9309 8919 9367 8925
rect 9861 8925 9873 8928
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8925 10195 8959
rect 10137 8919 10195 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 10321 8919 10379 8925
rect 10152 8888 10180 8919
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 12253 8959 12311 8965
rect 12253 8956 12265 8959
rect 11204 8928 12265 8956
rect 11204 8916 11210 8928
rect 12253 8925 12265 8928
rect 12299 8925 12311 8959
rect 12253 8919 12311 8925
rect 12526 8916 12532 8968
rect 12584 8916 12590 8968
rect 12618 8916 12624 8968
rect 12676 8916 12682 8968
rect 13078 8916 13084 8968
rect 13136 8956 13142 8968
rect 13173 8959 13231 8965
rect 13173 8956 13185 8959
rect 13136 8928 13185 8956
rect 13136 8916 13142 8928
rect 13173 8925 13185 8928
rect 13219 8925 13231 8959
rect 13173 8919 13231 8925
rect 9048 8860 10180 8888
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 12713 8891 12771 8897
rect 12713 8888 12725 8891
rect 12032 8860 12725 8888
rect 12032 8848 12038 8860
rect 12713 8857 12725 8860
rect 12759 8857 12771 8891
rect 12713 8851 12771 8857
rect 6880 8792 7328 8820
rect 6880 8780 6886 8792
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8481 8823 8539 8829
rect 8481 8820 8493 8823
rect 8168 8792 8493 8820
rect 8168 8780 8174 8792
rect 8481 8789 8493 8792
rect 8527 8789 8539 8823
rect 8481 8783 8539 8789
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 9398 8820 9404 8832
rect 8619 8792 9404 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 12066 8780 12072 8832
rect 12124 8780 12130 8832
rect 12434 8780 12440 8832
rect 12492 8780 12498 8832
rect 13354 8780 13360 8832
rect 13412 8780 13418 8832
rect 1104 8730 13800 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 13800 8730
rect 1104 8656 13800 8678
rect 1670 8576 1676 8628
rect 1728 8616 1734 8628
rect 2501 8619 2559 8625
rect 2501 8616 2513 8619
rect 1728 8588 2513 8616
rect 1728 8576 1734 8588
rect 2501 8585 2513 8588
rect 2547 8585 2559 8619
rect 2501 8579 2559 8585
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2648 8588 2973 8616
rect 2648 8576 2654 8588
rect 2961 8585 2973 8588
rect 3007 8616 3019 8619
rect 5626 8616 5632 8628
rect 3007 8588 5632 8616
rect 3007 8585 3019 8588
rect 2961 8579 3019 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 6086 8576 6092 8628
rect 6144 8616 6150 8628
rect 6181 8619 6239 8625
rect 6181 8616 6193 8619
rect 6144 8588 6193 8616
rect 6144 8576 6150 8588
rect 6181 8585 6193 8588
rect 6227 8585 6239 8619
rect 6546 8616 6552 8628
rect 6181 8579 6239 8585
rect 6288 8588 6552 8616
rect 2225 8551 2283 8557
rect 2225 8517 2237 8551
rect 2271 8548 2283 8551
rect 2406 8548 2412 8560
rect 2271 8520 2412 8548
rect 2271 8517 2283 8520
rect 2225 8511 2283 8517
rect 2406 8508 2412 8520
rect 2464 8548 2470 8560
rect 3881 8551 3939 8557
rect 3881 8548 3893 8551
rect 2464 8520 3893 8548
rect 2464 8508 2470 8520
rect 3881 8517 3893 8520
rect 3927 8548 3939 8551
rect 6288 8548 6316 8588
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 7006 8616 7012 8628
rect 6687 8588 7012 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 8294 8616 8300 8628
rect 7116 8588 8300 8616
rect 3927 8520 4016 8548
rect 3927 8517 3939 8520
rect 3881 8511 3939 8517
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 2866 8480 2872 8492
rect 1820 8452 2872 8480
rect 1820 8440 1826 8452
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 3988 8489 4016 8520
rect 4172 8520 6316 8548
rect 4172 8489 4200 8520
rect 6362 8508 6368 8560
rect 6420 8508 6426 8560
rect 3973 8483 4031 8489
rect 3973 8449 3985 8483
rect 4019 8449 4031 8483
rect 3973 8443 4031 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 2774 8304 2780 8356
rect 2832 8344 2838 8356
rect 3068 8344 3096 8375
rect 3326 8372 3332 8424
rect 3384 8372 3390 8424
rect 2832 8316 3096 8344
rect 2832 8304 2838 8316
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4172 8344 4200 8443
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5813 8483 5871 8489
rect 5813 8480 5825 8483
rect 5776 8452 5825 8480
rect 5776 8440 5782 8452
rect 5813 8449 5825 8452
rect 5859 8449 5871 8483
rect 5813 8443 5871 8449
rect 6454 8440 6460 8492
rect 6512 8480 6518 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6512 8452 6561 8480
rect 6512 8440 6518 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6638 8440 6644 8492
rect 6696 8480 6702 8492
rect 7116 8480 7144 8588
rect 8294 8576 8300 8588
rect 8352 8576 8358 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8996 8588 9045 8616
rect 8996 8576 9002 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9033 8579 9091 8585
rect 9122 8576 9128 8628
rect 9180 8576 9186 8628
rect 11333 8619 11391 8625
rect 11333 8585 11345 8619
rect 11379 8616 11391 8619
rect 12618 8616 12624 8628
rect 11379 8588 12624 8616
rect 11379 8585 11391 8588
rect 11333 8579 11391 8585
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 8202 8508 8208 8560
rect 8260 8548 8266 8560
rect 10965 8551 11023 8557
rect 8260 8520 9260 8548
rect 8260 8508 8266 8520
rect 6696 8452 7144 8480
rect 6696 8440 6702 8452
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 8297 8483 8355 8489
rect 8297 8480 8309 8483
rect 8168 8452 8309 8480
rect 8168 8440 8174 8452
rect 8297 8449 8309 8452
rect 8343 8449 8355 8483
rect 8297 8443 8355 8449
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 9133 8483 9191 8489
rect 9133 8449 9145 8483
rect 9179 8480 9191 8483
rect 9232 8480 9260 8520
rect 10965 8517 10977 8551
rect 11011 8548 11023 8551
rect 11054 8548 11060 8560
rect 11011 8520 11060 8548
rect 11011 8517 11023 8520
rect 10965 8511 11023 8517
rect 11054 8508 11060 8520
rect 11112 8508 11118 8560
rect 11181 8551 11239 8557
rect 11181 8517 11193 8551
rect 11227 8548 11239 8551
rect 11882 8548 11888 8560
rect 11227 8520 11888 8548
rect 11227 8517 11239 8520
rect 11181 8511 11239 8517
rect 11882 8508 11888 8520
rect 11940 8508 11946 8560
rect 12802 8508 12808 8560
rect 12860 8508 12866 8560
rect 9179 8452 9260 8480
rect 9309 8483 9367 8489
rect 9179 8449 9191 8452
rect 9133 8443 9191 8449
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9398 8480 9404 8492
rect 9355 8452 9404 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 5350 8372 5356 8424
rect 5408 8412 5414 8424
rect 5905 8415 5963 8421
rect 5905 8412 5917 8415
rect 5408 8384 5917 8412
rect 5408 8372 5414 8384
rect 5905 8381 5917 8384
rect 5951 8412 5963 8415
rect 8202 8412 8208 8424
rect 5951 8384 8208 8412
rect 5951 8381 5963 8384
rect 5905 8375 5963 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 3752 8316 4200 8344
rect 3752 8304 3758 8316
rect 4522 8304 4528 8356
rect 4580 8344 4586 8356
rect 5810 8344 5816 8356
rect 4580 8316 5816 8344
rect 4580 8304 4586 8316
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6178 8304 6184 8356
rect 6236 8344 6242 8356
rect 8404 8344 8432 8375
rect 8570 8372 8576 8424
rect 8628 8412 8634 8424
rect 9033 8415 9091 8421
rect 9033 8412 9045 8415
rect 8628 8384 9045 8412
rect 8628 8372 8634 8384
rect 9033 8381 9045 8384
rect 9079 8381 9091 8415
rect 9033 8375 9091 8381
rect 9214 8372 9220 8424
rect 9272 8412 9278 8424
rect 11238 8412 11244 8424
rect 9272 8384 11244 8412
rect 9272 8372 9278 8384
rect 11238 8372 11244 8384
rect 11296 8372 11302 8424
rect 11422 8372 11428 8424
rect 11480 8412 11486 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 11480 8384 11529 8412
rect 11480 8372 11486 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 11790 8372 11796 8424
rect 11848 8372 11854 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12526 8412 12532 8424
rect 11940 8384 12532 8412
rect 11940 8372 11946 8384
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 6236 8316 8984 8344
rect 6236 8304 6242 8316
rect 4062 8236 4068 8288
rect 4120 8236 4126 8288
rect 5074 8236 5080 8288
rect 5132 8276 5138 8288
rect 5626 8276 5632 8288
rect 5132 8248 5632 8276
rect 5132 8236 5138 8248
rect 5626 8236 5632 8248
rect 5684 8276 5690 8288
rect 5997 8279 6055 8285
rect 5997 8276 6009 8279
rect 5684 8248 6009 8276
rect 5684 8236 5690 8248
rect 5997 8245 6009 8248
rect 6043 8276 6055 8279
rect 6730 8276 6736 8288
rect 6043 8248 6736 8276
rect 6043 8245 6055 8248
rect 5997 8239 6055 8245
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 8662 8236 8668 8288
rect 8720 8236 8726 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 8849 8279 8907 8285
rect 8849 8276 8861 8279
rect 8812 8248 8861 8276
rect 8812 8236 8818 8248
rect 8849 8245 8861 8248
rect 8895 8245 8907 8279
rect 8956 8276 8984 8316
rect 9646 8316 11192 8344
rect 9646 8276 9674 8316
rect 11164 8288 11192 8316
rect 8956 8248 9674 8276
rect 8849 8239 8907 8245
rect 11146 8236 11152 8288
rect 11204 8236 11210 8288
rect 13262 8236 13268 8288
rect 13320 8236 13326 8288
rect 1104 8186 13800 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 13800 8186
rect 1104 8112 13800 8134
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 2746 8044 4445 8072
rect 2746 8004 2774 8044
rect 4433 8041 4445 8044
rect 4479 8041 4491 8075
rect 4433 8035 4491 8041
rect 5074 8032 5080 8084
rect 5132 8032 5138 8084
rect 5350 8032 5356 8084
rect 5408 8072 5414 8084
rect 5718 8072 5724 8084
rect 5408 8044 5724 8072
rect 5408 8032 5414 8044
rect 5718 8032 5724 8044
rect 5776 8072 5782 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5776 8044 5917 8072
rect 5776 8032 5782 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 5905 8035 5963 8041
rect 11146 8032 11152 8084
rect 11204 8032 11210 8084
rect 11790 8032 11796 8084
rect 11848 8072 11854 8084
rect 12253 8075 12311 8081
rect 12253 8072 12265 8075
rect 11848 8044 12265 8072
rect 11848 8032 11854 8044
rect 12253 8041 12265 8044
rect 12299 8041 12311 8075
rect 12253 8035 12311 8041
rect 13354 8032 13360 8084
rect 13412 8032 13418 8084
rect 5092 8004 5120 8032
rect 2424 7976 2774 8004
rect 5000 7976 5120 8004
rect 5445 8007 5503 8013
rect 2038 7828 2044 7880
rect 2096 7828 2102 7880
rect 2130 7828 2136 7880
rect 2188 7828 2194 7880
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2424 7868 2452 7976
rect 3326 7936 3332 7948
rect 2516 7908 3332 7936
rect 2516 7877 2544 7908
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 3786 7896 3792 7948
rect 3844 7896 3850 7948
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 4430 7936 4436 7948
rect 4295 7908 4436 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 4430 7896 4436 7908
rect 4488 7896 4494 7948
rect 4614 7896 4620 7948
rect 4672 7896 4678 7948
rect 2363 7840 2452 7868
rect 2501 7871 2559 7877
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 2501 7837 2513 7871
rect 2547 7837 2559 7871
rect 2501 7831 2559 7837
rect 2590 7828 2596 7880
rect 2648 7868 2654 7880
rect 2777 7871 2835 7877
rect 2777 7868 2789 7871
rect 2648 7840 2789 7868
rect 2648 7828 2654 7840
rect 2777 7837 2789 7840
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7870 4215 7871
rect 4203 7868 4292 7870
rect 4632 7868 4660 7896
rect 4203 7842 4660 7868
rect 4203 7837 4215 7842
rect 4264 7840 4660 7842
rect 4801 7871 4859 7877
rect 4157 7831 4215 7837
rect 4801 7837 4813 7871
rect 4847 7868 4859 7871
rect 5000 7868 5028 7976
rect 5445 7973 5457 8007
rect 5491 8004 5503 8007
rect 6454 8004 6460 8016
rect 5491 7976 6460 8004
rect 5491 7973 5503 7976
rect 5445 7967 5503 7973
rect 6454 7964 6460 7976
rect 6512 7964 6518 8016
rect 8846 7964 8852 8016
rect 8904 8004 8910 8016
rect 11425 8007 11483 8013
rect 11425 8004 11437 8007
rect 8904 7976 11437 8004
rect 8904 7964 8910 7976
rect 11425 7973 11437 7976
rect 11471 7973 11483 8007
rect 11425 7967 11483 7973
rect 5077 7939 5135 7945
rect 5077 7905 5089 7939
rect 5123 7936 5135 7939
rect 5626 7936 5632 7948
rect 5123 7908 5632 7936
rect 5123 7905 5135 7908
rect 5077 7899 5135 7905
rect 5626 7896 5632 7908
rect 5684 7936 5690 7948
rect 5813 7939 5871 7945
rect 5813 7936 5825 7939
rect 5684 7908 5825 7936
rect 5684 7896 5690 7908
rect 5813 7905 5825 7908
rect 5859 7936 5871 7939
rect 6086 7936 6092 7948
rect 5859 7908 6092 7936
rect 5859 7905 5871 7908
rect 5813 7899 5871 7905
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 6641 7939 6699 7945
rect 6641 7936 6653 7939
rect 6319 7908 6653 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 6641 7905 6653 7908
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 11149 7939 11207 7945
rect 11149 7936 11161 7939
rect 11112 7908 11161 7936
rect 11112 7896 11118 7908
rect 11149 7905 11161 7908
rect 11195 7936 11207 7939
rect 11195 7908 12480 7936
rect 11195 7905 11207 7908
rect 11149 7899 11207 7905
rect 4847 7840 5028 7868
rect 5261 7871 5319 7877
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 5261 7837 5273 7871
rect 5307 7868 5319 7871
rect 5442 7868 5448 7880
rect 5307 7840 5448 7868
rect 5307 7837 5319 7840
rect 5261 7831 5319 7837
rect 5442 7828 5448 7840
rect 5500 7828 5506 7880
rect 5534 7828 5540 7880
rect 5592 7828 5598 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 5997 7871 6055 7877
rect 5997 7837 6009 7871
rect 6043 7868 6055 7871
rect 6546 7868 6552 7880
rect 6043 7840 6552 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 2409 7803 2467 7809
rect 2409 7769 2421 7803
rect 2455 7800 2467 7803
rect 4062 7800 4068 7812
rect 2455 7772 4068 7800
rect 2455 7769 2467 7772
rect 2409 7763 2467 7769
rect 4062 7760 4068 7772
rect 4120 7760 4126 7812
rect 4617 7803 4675 7809
rect 4617 7769 4629 7803
rect 4663 7800 4675 7803
rect 4706 7800 4712 7812
rect 4663 7772 4712 7800
rect 4663 7769 4675 7772
rect 4617 7763 4675 7769
rect 4706 7760 4712 7772
rect 4764 7760 4770 7812
rect 4985 7803 5043 7809
rect 4985 7769 4997 7803
rect 5031 7800 5043 7803
rect 5350 7800 5356 7812
rect 5031 7772 5356 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 5350 7760 5356 7772
rect 5408 7760 5414 7812
rect 5736 7800 5764 7831
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7868 6791 7871
rect 8570 7868 8576 7880
rect 6779 7840 8576 7868
rect 6779 7837 6791 7840
rect 6733 7831 6791 7837
rect 8570 7828 8576 7840
rect 8628 7828 8634 7880
rect 9214 7828 9220 7880
rect 9272 7828 9278 7880
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9582 7868 9588 7880
rect 9447 7840 9588 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 11238 7828 11244 7880
rect 11296 7828 11302 7880
rect 11532 7877 11560 7908
rect 12452 7880 12480 7908
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 6822 7800 6828 7812
rect 5736 7772 6828 7800
rect 1581 7735 1639 7741
rect 1581 7701 1593 7735
rect 1627 7732 1639 7735
rect 1854 7732 1860 7744
rect 1627 7704 1860 7732
rect 1627 7701 1639 7704
rect 1581 7695 1639 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2682 7692 2688 7744
rect 2740 7692 2746 7744
rect 3326 7692 3332 7744
rect 3384 7692 3390 7744
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 5736 7732 5764 7772
rect 6822 7760 6828 7772
rect 6880 7760 6886 7812
rect 11146 7760 11152 7812
rect 11204 7800 11210 7812
rect 11624 7800 11652 7831
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 11974 7828 11980 7880
rect 12032 7828 12038 7880
rect 12066 7828 12072 7880
rect 12124 7828 12130 7880
rect 12250 7868 12256 7880
rect 12176 7840 12256 7868
rect 11204 7772 11652 7800
rect 11204 7760 11210 7772
rect 4948 7704 5764 7732
rect 4948 7692 4954 7704
rect 6362 7692 6368 7744
rect 6420 7692 6426 7744
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 9490 7732 9496 7744
rect 9447 7704 9496 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 9490 7692 9496 7704
rect 9548 7692 9554 7744
rect 10873 7735 10931 7741
rect 10873 7701 10885 7735
rect 10919 7732 10931 7735
rect 11054 7732 11060 7744
rect 10919 7704 11060 7732
rect 10919 7701 10931 7704
rect 10873 7695 10931 7701
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11624 7732 11652 7772
rect 11767 7803 11825 7809
rect 11767 7769 11779 7803
rect 11813 7800 11825 7803
rect 12176 7800 12204 7840
rect 12250 7828 12256 7840
rect 12308 7828 12314 7880
rect 12434 7828 12440 7880
rect 12492 7868 12498 7880
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12492 7840 12541 7868
rect 12492 7828 12498 7840
rect 12529 7837 12541 7840
rect 12575 7868 12587 7871
rect 12802 7868 12808 7880
rect 12575 7840 12808 7868
rect 12575 7837 12587 7840
rect 12529 7831 12587 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 13173 7871 13231 7877
rect 13173 7868 13185 7871
rect 12912 7840 13185 7868
rect 11813 7772 12204 7800
rect 12268 7772 12572 7800
rect 11813 7769 11825 7772
rect 11767 7763 11825 7769
rect 12268 7732 12296 7772
rect 11624 7704 12296 7732
rect 12342 7692 12348 7744
rect 12400 7692 12406 7744
rect 12544 7732 12572 7772
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 12713 7803 12771 7809
rect 12713 7800 12725 7803
rect 12676 7772 12725 7800
rect 12676 7760 12682 7772
rect 12713 7769 12725 7772
rect 12759 7769 12771 7803
rect 12713 7763 12771 7769
rect 12912 7732 12940 7840
rect 13173 7837 13185 7840
rect 13219 7868 13231 7871
rect 13262 7868 13268 7880
rect 13219 7840 13268 7868
rect 13219 7837 13231 7840
rect 13173 7831 13231 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 12544 7704 12940 7732
rect 12986 7692 12992 7744
rect 13044 7692 13050 7744
rect 1104 7642 13800 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 13800 7642
rect 1104 7568 13800 7590
rect 1673 7531 1731 7537
rect 1673 7497 1685 7531
rect 1719 7528 1731 7531
rect 2498 7528 2504 7540
rect 1719 7500 2504 7528
rect 1719 7497 1731 7500
rect 1673 7491 1731 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 2590 7488 2596 7540
rect 2648 7488 2654 7540
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6227 7500 6561 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 6914 7488 6920 7540
rect 6972 7488 6978 7540
rect 8754 7488 8760 7540
rect 8812 7528 8818 7540
rect 8812 7500 9168 7528
rect 8812 7488 8818 7500
rect 2038 7420 2044 7472
rect 2096 7460 2102 7472
rect 2608 7460 2636 7488
rect 2961 7463 3019 7469
rect 2961 7460 2973 7463
rect 2096 7432 2973 7460
rect 2096 7420 2102 7432
rect 2961 7429 2973 7432
rect 3007 7429 3019 7463
rect 2961 7423 3019 7429
rect 3513 7463 3571 7469
rect 3513 7429 3525 7463
rect 3559 7460 3571 7463
rect 3878 7460 3884 7472
rect 3559 7432 3884 7460
rect 3559 7429 3571 7432
rect 3513 7423 3571 7429
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 4341 7463 4399 7469
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 5258 7460 5264 7472
rect 4387 7432 5264 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 5258 7420 5264 7432
rect 5316 7420 5322 7472
rect 6362 7420 6368 7472
rect 6420 7420 6426 7472
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 9033 7463 9091 7469
rect 9033 7460 9045 7463
rect 6880 7432 9045 7460
rect 6880 7420 6886 7432
rect 9033 7429 9045 7432
rect 9079 7429 9091 7463
rect 9140 7460 9168 7500
rect 9214 7488 9220 7540
rect 9272 7488 9278 7540
rect 9306 7488 9312 7540
rect 9364 7488 9370 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10594 7528 10600 7540
rect 9999 7500 10600 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 12802 7488 12808 7540
rect 12860 7528 12866 7540
rect 13357 7531 13415 7537
rect 13357 7528 13369 7531
rect 12860 7500 13369 7528
rect 12860 7488 12866 7500
rect 13357 7497 13369 7500
rect 13403 7497 13415 7531
rect 13357 7491 13415 7497
rect 9324 7460 9352 7488
rect 9140 7432 9444 7460
rect 9033 7423 9091 7429
rect 1670 7352 1676 7404
rect 1728 7352 1734 7404
rect 1854 7352 1860 7404
rect 1912 7352 1918 7404
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7392 2467 7395
rect 2455 7364 2544 7392
rect 2455 7361 2467 7364
rect 2409 7355 2467 7361
rect 2516 7256 2544 7364
rect 2590 7352 2596 7404
rect 2648 7352 2654 7404
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3602 7352 3608 7404
rect 3660 7352 3666 7404
rect 3786 7401 3792 7404
rect 3752 7395 3792 7401
rect 3752 7361 3764 7395
rect 3752 7355 3792 7361
rect 3786 7352 3792 7355
rect 3844 7352 3850 7404
rect 4430 7352 4436 7404
rect 4488 7392 4494 7404
rect 5169 7395 5227 7401
rect 5169 7392 5181 7395
rect 4488 7364 5181 7392
rect 4488 7352 4494 7364
rect 5169 7361 5181 7364
rect 5215 7392 5227 7395
rect 5442 7392 5448 7404
rect 5215 7364 5448 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 2682 7284 2688 7336
rect 2740 7324 2746 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 2740 7296 3985 7324
rect 2740 7284 2746 7296
rect 3973 7293 3985 7296
rect 4019 7293 4031 7327
rect 3973 7287 4031 7293
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 5350 7324 5356 7336
rect 5307 7296 5356 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 5350 7284 5356 7296
rect 5408 7284 5414 7336
rect 5537 7327 5595 7333
rect 5537 7293 5549 7327
rect 5583 7324 5595 7327
rect 5721 7327 5779 7333
rect 5721 7324 5733 7327
rect 5583 7296 5733 7324
rect 5583 7293 5595 7296
rect 5537 7287 5595 7293
rect 5721 7293 5733 7296
rect 5767 7293 5779 7327
rect 5828 7324 5856 7355
rect 6178 7352 6184 7404
rect 6236 7392 6242 7404
rect 6641 7395 6699 7401
rect 6641 7392 6653 7395
rect 6236 7364 6653 7392
rect 6236 7352 6242 7364
rect 6641 7361 6653 7364
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 7098 7392 7104 7404
rect 6779 7364 7104 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 7098 7352 7104 7364
rect 7156 7352 7162 7404
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 8846 7324 8852 7336
rect 5828 7296 8852 7324
rect 5721 7287 5779 7293
rect 8846 7284 8852 7296
rect 8904 7324 8910 7336
rect 8956 7324 8984 7355
rect 9122 7352 9128 7404
rect 9180 7352 9186 7404
rect 9306 7352 9312 7404
rect 9364 7352 9370 7404
rect 9416 7401 9444 7432
rect 9490 7420 9496 7472
rect 9548 7420 9554 7472
rect 12894 7420 12900 7472
rect 12952 7420 12958 7472
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 9766 7352 9772 7404
rect 9824 7352 9830 7404
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 10045 7395 10103 7401
rect 10045 7392 10057 7395
rect 9916 7364 10057 7392
rect 9916 7352 9922 7364
rect 10045 7361 10057 7364
rect 10091 7361 10103 7395
rect 10045 7355 10103 7361
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 8904 7296 8984 7324
rect 9677 7327 9735 7333
rect 8904 7284 8910 7296
rect 9677 7293 9689 7327
rect 9723 7324 9735 7327
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 9723 7296 10149 7324
rect 9723 7293 9735 7296
rect 9677 7287 9735 7293
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 11422 7284 11428 7336
rect 11480 7324 11486 7336
rect 11609 7327 11667 7333
rect 11609 7324 11621 7327
rect 11480 7296 11621 7324
rect 11480 7284 11486 7296
rect 11609 7293 11621 7296
rect 11655 7293 11667 7327
rect 11609 7287 11667 7293
rect 11882 7284 11888 7336
rect 11940 7284 11946 7336
rect 2958 7256 2964 7268
rect 2516 7228 2964 7256
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3881 7191 3939 7197
rect 3881 7188 3893 7191
rect 3292 7160 3893 7188
rect 3292 7148 3298 7160
rect 3881 7157 3893 7160
rect 3927 7157 3939 7191
rect 3881 7151 3939 7157
rect 9490 7148 9496 7200
rect 9548 7148 9554 7200
rect 1104 7098 13800 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 13800 7098
rect 1104 7024 13800 7046
rect 3602 6944 3608 6996
rect 3660 6984 3666 6996
rect 4433 6987 4491 6993
rect 4433 6984 4445 6987
rect 3660 6956 4445 6984
rect 3660 6944 3666 6956
rect 4433 6953 4445 6956
rect 4479 6953 4491 6987
rect 4433 6947 4491 6953
rect 11793 6987 11851 6993
rect 11793 6953 11805 6987
rect 11839 6984 11851 6987
rect 11882 6984 11888 6996
rect 11839 6956 11888 6984
rect 11839 6953 11851 6956
rect 11793 6947 11851 6953
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 3142 6916 3148 6928
rect 2976 6888 3148 6916
rect 2038 6808 2044 6860
rect 2096 6808 2102 6860
rect 2976 6857 3004 6888
rect 3142 6876 3148 6888
rect 3200 6916 3206 6928
rect 3200 6888 3556 6916
rect 3200 6876 3206 6888
rect 2961 6851 3019 6857
rect 2961 6817 2973 6851
rect 3007 6817 3019 6851
rect 2961 6811 3019 6817
rect 3050 6808 3056 6860
rect 3108 6808 3114 6860
rect 3528 6848 3556 6888
rect 8846 6876 8852 6928
rect 8904 6916 8910 6928
rect 9585 6919 9643 6925
rect 9585 6916 9597 6919
rect 8904 6888 9597 6916
rect 8904 6876 8910 6888
rect 9585 6885 9597 6888
rect 9631 6916 9643 6919
rect 10226 6916 10232 6928
rect 9631 6888 10232 6916
rect 9631 6885 9643 6888
rect 9585 6879 9643 6885
rect 10226 6876 10232 6888
rect 10284 6916 10290 6928
rect 10284 6888 10640 6916
rect 10284 6876 10290 6888
rect 4338 6848 4344 6860
rect 3528 6820 4344 6848
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 3068 6712 3096 6808
rect 3326 6740 3332 6792
rect 3384 6740 3390 6792
rect 3528 6789 3556 6820
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 8478 6808 8484 6860
rect 8536 6808 8542 6860
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6817 8815 6851
rect 8757 6811 8815 6817
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6848 8999 6851
rect 9030 6848 9036 6860
rect 8987 6820 9036 6848
rect 8987 6817 8999 6820
rect 8941 6811 8999 6817
rect 3513 6783 3571 6789
rect 3513 6749 3525 6783
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3786 6740 3792 6792
rect 3844 6740 3850 6792
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4254 6783 4312 6789
rect 3936 6752 3981 6780
rect 3936 6740 3942 6752
rect 4254 6749 4266 6783
rect 4300 6749 4312 6783
rect 4254 6743 4312 6749
rect 3142 6712 3148 6724
rect 3068 6684 3148 6712
rect 3142 6672 3148 6684
rect 3200 6672 3206 6724
rect 2498 6604 2504 6656
rect 2556 6604 2562 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3344 6644 3372 6740
rect 3421 6715 3479 6721
rect 3421 6681 3433 6715
rect 3467 6712 3479 6715
rect 4065 6715 4123 6721
rect 4065 6712 4077 6715
rect 3467 6684 4077 6712
rect 3467 6681 3479 6684
rect 3421 6675 3479 6681
rect 4065 6681 4077 6684
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 4154 6672 4160 6724
rect 4212 6672 4218 6724
rect 2915 6616 3372 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 4264 6644 4292 6743
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8389 6783 8447 6789
rect 8389 6780 8401 6783
rect 8260 6752 8401 6780
rect 8260 6740 8266 6752
rect 8389 6749 8401 6752
rect 8435 6749 8447 6783
rect 8772 6780 8800 6811
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 9766 6848 9772 6860
rect 9140 6820 9772 6848
rect 9140 6780 9168 6820
rect 9766 6808 9772 6820
rect 9824 6848 9830 6860
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 9824 6820 10057 6848
rect 9824 6808 9830 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 8772 6752 9168 6780
rect 8389 6743 8447 6749
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9732 6752 10088 6780
rect 9732 6740 9738 6752
rect 9309 6715 9367 6721
rect 9309 6681 9321 6715
rect 9355 6712 9367 6715
rect 10060 6712 10088 6752
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10612 6789 10640 6888
rect 12342 6848 12348 6860
rect 11992 6820 12348 6848
rect 11992 6789 12020 6820
rect 12342 6808 12348 6820
rect 12400 6808 12406 6860
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12492 6820 12756 6848
rect 12492 6808 12498 6820
rect 10413 6783 10471 6789
rect 10413 6749 10425 6783
rect 10459 6749 10471 6783
rect 10413 6743 10471 6749
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 11977 6743 12035 6749
rect 12452 6752 12541 6780
rect 10428 6712 10456 6743
rect 12452 6724 12480 6752
rect 12529 6749 12541 6752
rect 12575 6780 12587 6783
rect 12618 6780 12624 6792
rect 12575 6752 12624 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 12618 6740 12624 6752
rect 12676 6740 12682 6792
rect 12728 6789 12756 6820
rect 12713 6783 12771 6789
rect 12713 6749 12725 6783
rect 12759 6749 12771 6783
rect 12713 6743 12771 6749
rect 9355 6684 9812 6712
rect 10060 6684 10456 6712
rect 12069 6715 12127 6721
rect 9355 6681 9367 6684
rect 9309 6675 9367 6681
rect 3660 6616 4292 6644
rect 3660 6604 3666 6616
rect 9398 6604 9404 6656
rect 9456 6604 9462 6656
rect 9784 6653 9812 6684
rect 12069 6681 12081 6715
rect 12115 6681 12127 6715
rect 12069 6675 12127 6681
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6613 9827 6647
rect 9769 6607 9827 6613
rect 10410 6604 10416 6656
rect 10468 6604 10474 6656
rect 12084 6644 12112 6675
rect 12158 6672 12164 6724
rect 12216 6672 12222 6724
rect 12250 6672 12256 6724
rect 12308 6721 12314 6724
rect 12308 6715 12337 6721
rect 12325 6681 12337 6715
rect 12308 6675 12337 6681
rect 12308 6672 12314 6675
rect 12434 6672 12440 6724
rect 12492 6672 12498 6724
rect 12621 6647 12679 6653
rect 12621 6644 12633 6647
rect 12084 6616 12633 6644
rect 12621 6613 12633 6616
rect 12667 6613 12679 6647
rect 12621 6607 12679 6613
rect 1104 6554 13800 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 13800 6554
rect 1104 6480 13800 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 2866 6440 2872 6452
rect 1627 6412 2872 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 1670 6332 1676 6384
rect 1728 6332 1734 6384
rect 2424 6381 2452 6412
rect 2866 6400 2872 6412
rect 2924 6440 2930 6452
rect 4249 6443 4307 6449
rect 2924 6412 4108 6440
rect 2924 6400 2930 6412
rect 2409 6375 2467 6381
rect 2409 6341 2421 6375
rect 2455 6341 2467 6375
rect 2409 6335 2467 6341
rect 2498 6332 2504 6384
rect 2556 6372 2562 6384
rect 2777 6375 2835 6381
rect 2777 6372 2789 6375
rect 2556 6344 2789 6372
rect 2556 6332 2562 6344
rect 2777 6341 2789 6344
rect 2823 6341 2835 6375
rect 2777 6335 2835 6341
rect 934 6264 940 6316
rect 992 6304 998 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 992 6276 1409 6304
rect 992 6264 998 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 4080 6304 4108 6412
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 4338 6440 4344 6452
rect 4295 6412 4344 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4338 6400 4344 6412
rect 4396 6440 4402 6452
rect 5169 6443 5227 6449
rect 4396 6412 5120 6440
rect 4396 6400 4402 6412
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 4433 6375 4491 6381
rect 4433 6372 4445 6375
rect 4212 6344 4445 6372
rect 4212 6332 4218 6344
rect 4433 6341 4445 6344
rect 4479 6341 4491 6375
rect 5092 6372 5120 6412
rect 5169 6409 5181 6443
rect 5215 6440 5227 6443
rect 5350 6440 5356 6452
rect 5215 6412 5356 6440
rect 5215 6409 5227 6412
rect 5169 6403 5227 6409
rect 5350 6400 5356 6412
rect 5408 6400 5414 6452
rect 6822 6440 6828 6452
rect 5828 6412 6828 6440
rect 5828 6384 5856 6412
rect 6822 6400 6828 6412
rect 6880 6440 6886 6452
rect 6880 6412 7052 6440
rect 6880 6400 6886 6412
rect 5442 6372 5448 6384
rect 5092 6344 5448 6372
rect 4433 6335 4491 6341
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 5810 6372 5816 6384
rect 5552 6344 5816 6372
rect 4706 6304 4712 6316
rect 3910 6276 4016 6304
rect 4080 6276 4712 6304
rect 1397 6267 1455 6273
rect 3988 6248 4016 6276
rect 4706 6264 4712 6276
rect 4764 6264 4770 6316
rect 4798 6264 4804 6316
rect 4856 6264 4862 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6273 5043 6307
rect 4985 6267 5043 6273
rect 2038 6196 2044 6248
rect 2096 6196 2102 6248
rect 2406 6196 2412 6248
rect 2464 6236 2470 6248
rect 2501 6239 2559 6245
rect 2501 6236 2513 6239
rect 2464 6208 2513 6236
rect 2464 6196 2470 6208
rect 2501 6205 2513 6208
rect 2547 6205 2559 6239
rect 2501 6199 2559 6205
rect 3970 6196 3976 6248
rect 4028 6196 4034 6248
rect 5000 6236 5028 6267
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5552 6304 5580 6344
rect 5810 6332 5816 6344
rect 5868 6332 5874 6384
rect 7024 6372 7052 6412
rect 8938 6400 8944 6452
rect 8996 6400 9002 6452
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9398 6440 9404 6452
rect 9355 6412 9404 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 10686 6440 10692 6452
rect 10643 6412 10692 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 12250 6440 12256 6452
rect 10836 6412 12256 6440
rect 10836 6400 10842 6412
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 7561 6375 7619 6381
rect 7561 6372 7573 6375
rect 7024 6344 7573 6372
rect 7561 6341 7573 6344
rect 7607 6341 7619 6375
rect 7777 6375 7835 6381
rect 7777 6372 7789 6375
rect 7561 6335 7619 6341
rect 7668 6344 7789 6372
rect 5408 6276 5580 6304
rect 5629 6307 5687 6313
rect 5408 6264 5414 6276
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 5718 6304 5724 6316
rect 5675 6276 5724 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6454 6264 6460 6316
rect 6512 6264 6518 6316
rect 6641 6307 6699 6313
rect 6641 6273 6653 6307
rect 6687 6273 6699 6307
rect 6641 6267 6699 6273
rect 5442 6236 5448 6248
rect 5000 6208 5448 6236
rect 5442 6196 5448 6208
rect 5500 6196 5506 6248
rect 5534 6196 5540 6248
rect 5592 6196 5598 6248
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 6546 6236 6552 6248
rect 6411 6208 6552 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 6656 6236 6684 6267
rect 6730 6264 6736 6316
rect 6788 6264 6794 6316
rect 6825 6307 6883 6313
rect 6825 6273 6837 6307
rect 6871 6304 6883 6307
rect 6914 6304 6920 6316
rect 6871 6276 6920 6304
rect 6871 6273 6883 6276
rect 6825 6267 6883 6273
rect 6914 6264 6920 6276
rect 6972 6264 6978 6316
rect 7098 6264 7104 6316
rect 7156 6264 7162 6316
rect 7006 6236 7012 6248
rect 6656 6208 7012 6236
rect 7006 6196 7012 6208
rect 7064 6196 7070 6248
rect 4798 6168 4804 6180
rect 3804 6140 4804 6168
rect 2130 6060 2136 6112
rect 2188 6060 2194 6112
rect 2271 6103 2329 6109
rect 2271 6069 2283 6103
rect 2317 6100 2329 6103
rect 2498 6100 2504 6112
rect 2317 6072 2504 6100
rect 2317 6069 2329 6072
rect 2271 6063 2329 6069
rect 2498 6060 2504 6072
rect 2556 6100 2562 6112
rect 3804 6100 3832 6140
rect 4798 6128 4804 6140
rect 4856 6128 4862 6180
rect 5552 6168 5580 6196
rect 7668 6168 7696 6344
rect 7777 6341 7789 6344
rect 7823 6372 7835 6375
rect 7823 6344 8340 6372
rect 7823 6341 7835 6344
rect 7777 6335 7835 6341
rect 8312 6316 8340 6344
rect 8754 6332 8760 6384
rect 8812 6332 8818 6384
rect 9125 6375 9183 6381
rect 9125 6341 9137 6375
rect 9171 6372 9183 6375
rect 10410 6372 10416 6384
rect 9171 6344 10416 6372
rect 9171 6341 9183 6344
rect 9125 6335 9183 6341
rect 10410 6332 10416 6344
rect 10468 6332 10474 6384
rect 11054 6332 11060 6384
rect 11112 6332 11118 6384
rect 8110 6304 8116 6316
rect 5552 6140 7696 6168
rect 7760 6276 8116 6304
rect 2556 6072 3832 6100
rect 2556 6060 2562 6072
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 7760 6109 7788 6276
rect 8110 6264 8116 6276
rect 8168 6304 8174 6316
rect 8205 6307 8263 6313
rect 8205 6304 8217 6307
rect 8168 6276 8217 6304
rect 8168 6264 8174 6276
rect 8205 6273 8217 6276
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8386 6264 8392 6316
rect 8444 6264 8450 6316
rect 9030 6264 9036 6316
rect 9088 6264 9094 6316
rect 9769 6307 9827 6313
rect 9769 6304 9781 6307
rect 9140 6276 9781 6304
rect 8573 6239 8631 6245
rect 8573 6205 8585 6239
rect 8619 6236 8631 6239
rect 8619 6208 8892 6236
rect 8619 6205 8631 6208
rect 8573 6199 8631 6205
rect 8018 6128 8024 6180
rect 8076 6128 8082 6180
rect 8864 6168 8892 6208
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9140 6236 9168 6276
rect 9769 6273 9781 6276
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10318 6264 10324 6316
rect 10376 6304 10382 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10376 6276 10793 6304
rect 10376 6264 10382 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 10781 6267 10839 6273
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6304 12219 6307
rect 12434 6304 12440 6316
rect 12207 6276 12440 6304
rect 12207 6273 12219 6276
rect 12161 6267 12219 6273
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 8996 6208 9168 6236
rect 8996 6196 9002 6208
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9401 6239 9459 6245
rect 9401 6236 9413 6239
rect 9272 6208 9413 6236
rect 9272 6196 9278 6208
rect 9401 6205 9413 6208
rect 9447 6205 9459 6239
rect 9401 6199 9459 6205
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 9677 6239 9735 6245
rect 9677 6236 9689 6239
rect 9548 6208 9689 6236
rect 9548 6196 9554 6208
rect 9677 6205 9689 6208
rect 9723 6205 9735 6239
rect 9677 6199 9735 6205
rect 10870 6196 10876 6248
rect 10928 6196 10934 6248
rect 9582 6168 9588 6180
rect 8496 6140 8708 6168
rect 8864 6140 9588 6168
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 5592 6072 7757 6100
rect 5592 6060 5598 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8496 6100 8524 6140
rect 7975 6072 8524 6100
rect 8680 6100 8708 6140
rect 9582 6128 9588 6140
rect 9640 6168 9646 6180
rect 10134 6168 10140 6180
rect 9640 6140 10140 6168
rect 9640 6128 9646 6140
rect 10134 6128 10140 6140
rect 10192 6128 10198 6180
rect 9674 6100 9680 6112
rect 8680 6072 9680 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 10686 6060 10692 6112
rect 10744 6100 10750 6112
rect 10781 6103 10839 6109
rect 10781 6100 10793 6103
rect 10744 6072 10793 6100
rect 10744 6060 10750 6072
rect 10781 6069 10793 6072
rect 10827 6069 10839 6103
rect 10781 6063 10839 6069
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 12069 6103 12127 6109
rect 12069 6100 12081 6103
rect 11112 6072 12081 6100
rect 11112 6060 11118 6072
rect 12069 6069 12081 6072
rect 12115 6069 12127 6103
rect 12069 6063 12127 6069
rect 1104 6010 13800 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 13800 6010
rect 1104 5936 13800 5958
rect 3234 5856 3240 5908
rect 3292 5856 3298 5908
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 3602 5896 3608 5908
rect 3467 5868 3608 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 3602 5856 3608 5868
rect 3660 5856 3666 5908
rect 6365 5899 6423 5905
rect 5644 5868 6316 5896
rect 2225 5831 2283 5837
rect 2225 5797 2237 5831
rect 2271 5828 2283 5831
rect 3786 5828 3792 5840
rect 2271 5800 3792 5828
rect 2271 5797 2283 5800
rect 2225 5791 2283 5797
rect 3786 5788 3792 5800
rect 3844 5788 3850 5840
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2961 5763 3019 5769
rect 1995 5732 2268 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 2240 5704 2268 5732
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 3050 5760 3056 5772
rect 3007 5732 3056 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 3050 5720 3056 5732
rect 3108 5720 3114 5772
rect 842 5652 848 5704
rect 900 5692 906 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 900 5664 1409 5692
rect 900 5652 906 5664
rect 1397 5661 1409 5664
rect 1443 5661 1455 5695
rect 1397 5655 1455 5661
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5692 1915 5695
rect 2130 5692 2136 5704
rect 1903 5664 2136 5692
rect 1903 5661 1915 5664
rect 1857 5655 1915 5661
rect 1581 5559 1639 5565
rect 1581 5525 1593 5559
rect 1627 5556 1639 5559
rect 1872 5556 1900 5655
rect 2130 5652 2136 5664
rect 2188 5652 2194 5704
rect 2222 5652 2228 5704
rect 2280 5652 2286 5704
rect 2869 5695 2927 5701
rect 2869 5692 2881 5695
rect 2746 5664 2881 5692
rect 2038 5584 2044 5636
rect 2096 5624 2102 5636
rect 2746 5624 2774 5664
rect 2869 5661 2881 5664
rect 2915 5661 2927 5695
rect 2869 5655 2927 5661
rect 3329 5695 3387 5701
rect 3329 5661 3341 5695
rect 3375 5661 3387 5695
rect 3329 5655 3387 5661
rect 3513 5695 3571 5701
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 4798 5692 4804 5704
rect 3559 5664 4804 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 2096 5596 2774 5624
rect 2096 5584 2102 5596
rect 2958 5584 2964 5636
rect 3016 5624 3022 5636
rect 3344 5624 3372 5655
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5644 5692 5672 5868
rect 5718 5788 5724 5840
rect 5776 5828 5782 5840
rect 5776 5800 6132 5828
rect 5776 5788 5782 5800
rect 5902 5720 5908 5772
rect 5960 5720 5966 5772
rect 6104 5760 6132 5800
rect 6178 5788 6184 5840
rect 6236 5788 6242 5840
rect 6288 5828 6316 5868
rect 6365 5865 6377 5899
rect 6411 5896 6423 5899
rect 6730 5896 6736 5908
rect 6411 5868 6736 5896
rect 6411 5865 6423 5868
rect 6365 5859 6423 5865
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 8021 5899 8079 5905
rect 8021 5865 8033 5899
rect 8067 5896 8079 5899
rect 8938 5896 8944 5908
rect 8067 5868 8944 5896
rect 8067 5865 8079 5868
rect 8021 5859 8079 5865
rect 8938 5856 8944 5868
rect 8996 5856 9002 5908
rect 9306 5856 9312 5908
rect 9364 5856 9370 5908
rect 10597 5899 10655 5905
rect 10597 5865 10609 5899
rect 10643 5896 10655 5899
rect 12434 5896 12440 5908
rect 10643 5868 12440 5896
rect 10643 5865 10655 5868
rect 10597 5859 10655 5865
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 8202 5828 8208 5840
rect 6288 5800 8208 5828
rect 8202 5788 8208 5800
rect 8260 5828 8266 5840
rect 8757 5831 8815 5837
rect 8260 5800 8340 5828
rect 8260 5788 8266 5800
rect 8312 5769 8340 5800
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 8846 5828 8852 5840
rect 8803 5800 8852 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 8846 5788 8852 5800
rect 8904 5788 8910 5840
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 9493 5831 9551 5837
rect 9493 5828 9505 5831
rect 9180 5800 9505 5828
rect 9180 5788 9186 5800
rect 9493 5797 9505 5800
rect 9539 5797 9551 5831
rect 9493 5791 9551 5797
rect 8297 5763 8355 5769
rect 6104 5732 8248 5760
rect 5813 5695 5871 5701
rect 5813 5692 5825 5695
rect 5644 5664 5825 5692
rect 5813 5661 5825 5664
rect 5859 5661 5871 5695
rect 5813 5655 5871 5661
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5692 6607 5695
rect 6638 5692 6644 5704
rect 6595 5664 6644 5692
rect 6595 5661 6607 5664
rect 6549 5655 6607 5661
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 6822 5692 6828 5704
rect 6779 5664 6828 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 6822 5652 6828 5664
rect 6880 5692 6886 5704
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 6880 5664 7941 5692
rect 6880 5652 6886 5664
rect 7929 5661 7941 5664
rect 7975 5692 7987 5695
rect 8018 5692 8024 5704
rect 7975 5664 8024 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8110 5652 8116 5704
rect 8168 5652 8174 5704
rect 8220 5692 8248 5732
rect 8297 5729 8309 5763
rect 8343 5729 8355 5763
rect 8297 5723 8355 5729
rect 8478 5720 8484 5772
rect 8536 5760 8542 5772
rect 8536 5732 10456 5760
rect 8536 5720 8542 5732
rect 8386 5692 8392 5704
rect 8220 5664 8392 5692
rect 8386 5652 8392 5664
rect 8444 5652 8450 5704
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8904 5664 9137 5692
rect 8904 5652 8910 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 9125 5655 9183 5661
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9585 5695 9643 5701
rect 9585 5692 9597 5695
rect 9401 5655 9459 5661
rect 9508 5664 9597 5692
rect 5442 5624 5448 5636
rect 3016 5596 5448 5624
rect 3016 5584 3022 5596
rect 5442 5584 5448 5596
rect 5500 5584 5506 5636
rect 6656 5624 6684 5652
rect 8941 5627 8999 5633
rect 8941 5624 8953 5627
rect 6656 5596 8953 5624
rect 8941 5593 8953 5596
rect 8987 5624 8999 5627
rect 9214 5624 9220 5636
rect 8987 5596 9220 5624
rect 8987 5593 8999 5596
rect 8941 5587 8999 5593
rect 9214 5584 9220 5596
rect 9272 5584 9278 5636
rect 9416 5624 9444 5655
rect 9324 5596 9444 5624
rect 1627 5528 1900 5556
rect 1627 5525 1639 5528
rect 1581 5519 1639 5525
rect 4798 5516 4804 5568
rect 4856 5556 4862 5568
rect 5350 5556 5356 5568
rect 4856 5528 5356 5556
rect 4856 5516 4862 5528
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6641 5559 6699 5565
rect 6641 5556 6653 5559
rect 6604 5528 6653 5556
rect 6604 5516 6610 5528
rect 6641 5525 6653 5528
rect 6687 5525 6699 5559
rect 6641 5519 6699 5525
rect 8110 5516 8116 5568
rect 8168 5556 8174 5568
rect 9324 5556 9352 5596
rect 8168 5528 9352 5556
rect 8168 5516 8174 5528
rect 9398 5516 9404 5568
rect 9456 5556 9462 5568
rect 9508 5556 9536 5664
rect 9585 5661 9597 5664
rect 9631 5661 9643 5695
rect 9585 5655 9643 5661
rect 10318 5652 10324 5704
rect 10376 5652 10382 5704
rect 10428 5701 10456 5732
rect 11422 5720 11428 5772
rect 11480 5720 11486 5772
rect 10413 5695 10471 5701
rect 10413 5661 10425 5695
rect 10459 5692 10471 5695
rect 10686 5692 10692 5704
rect 10459 5664 10692 5692
rect 10459 5661 10471 5664
rect 10413 5655 10471 5661
rect 10686 5652 10692 5664
rect 10744 5652 10750 5704
rect 11054 5652 11060 5704
rect 11112 5652 11118 5704
rect 11146 5652 11152 5704
rect 11204 5652 11210 5704
rect 12802 5652 12808 5704
rect 12860 5652 12866 5704
rect 10042 5584 10048 5636
rect 10100 5584 10106 5636
rect 10152 5596 10732 5624
rect 9456 5528 9536 5556
rect 9456 5516 9462 5528
rect 9858 5516 9864 5568
rect 9916 5556 9922 5568
rect 10152 5556 10180 5596
rect 9916 5528 10180 5556
rect 9916 5516 9922 5528
rect 10226 5516 10232 5568
rect 10284 5516 10290 5568
rect 10704 5556 10732 5596
rect 10778 5584 10784 5636
rect 10836 5633 10842 5636
rect 10836 5627 10885 5633
rect 10836 5593 10839 5627
rect 10873 5593 10885 5627
rect 10836 5587 10885 5593
rect 10965 5627 11023 5633
rect 10965 5593 10977 5627
rect 11011 5593 11023 5627
rect 10965 5587 11023 5593
rect 11333 5627 11391 5633
rect 11333 5593 11345 5627
rect 11379 5624 11391 5627
rect 11701 5627 11759 5633
rect 11701 5624 11713 5627
rect 11379 5596 11713 5624
rect 11379 5593 11391 5596
rect 11333 5587 11391 5593
rect 11701 5593 11713 5596
rect 11747 5593 11759 5627
rect 11701 5587 11759 5593
rect 10836 5584 10842 5587
rect 10980 5556 11008 5587
rect 13446 5584 13452 5636
rect 13504 5584 13510 5636
rect 12066 5556 12072 5568
rect 10704 5528 12072 5556
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 1104 5466 13800 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 13800 5466
rect 1104 5392 13800 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 2038 5352 2044 5364
rect 1627 5324 2044 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 2130 5312 2136 5364
rect 2188 5312 2194 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 5537 5355 5595 5361
rect 3108 5324 4936 5352
rect 3108 5312 3114 5324
rect 2056 5284 2084 5312
rect 2961 5287 3019 5293
rect 2961 5284 2973 5287
rect 2056 5256 2973 5284
rect 2961 5253 2973 5256
rect 3007 5253 3019 5287
rect 2961 5247 3019 5253
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 4798 5176 4804 5228
rect 4856 5176 4862 5228
rect 4908 5225 4936 5324
rect 5537 5321 5549 5355
rect 5583 5321 5595 5355
rect 5537 5315 5595 5321
rect 5552 5284 5580 5315
rect 7006 5312 7012 5364
rect 7064 5312 7070 5364
rect 11146 5312 11152 5364
rect 11204 5352 11210 5364
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 11204 5324 11529 5352
rect 11204 5312 11210 5324
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 12802 5312 12808 5364
rect 12860 5312 12866 5364
rect 5994 5284 6000 5296
rect 5552 5256 6000 5284
rect 5994 5244 6000 5256
rect 6052 5284 6058 5296
rect 6454 5284 6460 5296
rect 6052 5256 6460 5284
rect 6052 5244 6058 5256
rect 6454 5244 6460 5256
rect 6512 5284 6518 5296
rect 6512 5256 6776 5284
rect 6512 5244 6518 5256
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 4893 5179 4951 5185
rect 5092 5188 5181 5216
rect 2222 5108 2228 5160
rect 2280 5108 2286 5160
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5117 2467 5151
rect 3142 5148 3148 5160
rect 2409 5111 2467 5117
rect 2746 5120 3148 5148
rect 2424 5080 2452 5111
rect 2746 5080 2774 5120
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 2424 5052 2774 5080
rect 4908 5080 4936 5179
rect 5092 5157 5120 5188
rect 5169 5185 5181 5188
rect 5215 5216 5227 5219
rect 5442 5216 5448 5228
rect 5215 5188 5448 5216
rect 5215 5185 5227 5188
rect 5169 5179 5227 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 5813 5219 5871 5225
rect 5813 5216 5825 5219
rect 5776 5188 5825 5216
rect 5776 5176 5782 5188
rect 5813 5185 5825 5188
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 6144 5188 6377 5216
rect 6144 5176 6150 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 6748 5225 6776 5256
rect 10686 5244 10692 5296
rect 10744 5284 10750 5296
rect 12897 5287 12955 5293
rect 10744 5256 12020 5284
rect 10744 5244 10750 5256
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6733 5219 6791 5225
rect 6733 5185 6745 5219
rect 6779 5185 6791 5219
rect 6733 5179 6791 5185
rect 5077 5151 5135 5157
rect 5077 5117 5089 5151
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 5350 5148 5356 5160
rect 5307 5120 5356 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 5350 5108 5356 5120
rect 5408 5108 5414 5160
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6270 5148 6276 5160
rect 6227 5120 6276 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 5534 5080 5540 5092
rect 4908 5052 5540 5080
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 1765 5015 1823 5021
rect 1765 5012 1777 5015
rect 1728 4984 1777 5012
rect 1728 4972 1734 4984
rect 1765 4981 1777 4984
rect 1811 4981 1823 5015
rect 1765 4975 1823 4981
rect 2590 4972 2596 5024
rect 2648 4972 2654 5024
rect 4982 4972 4988 5024
rect 5040 4972 5046 5024
rect 5184 5021 5212 5052
rect 5534 5040 5540 5052
rect 5592 5040 5598 5092
rect 5920 5080 5948 5111
rect 6270 5108 6276 5120
rect 6328 5148 6334 5160
rect 6656 5148 6684 5179
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 11992 5225 12020 5256
rect 12897 5253 12909 5287
rect 12943 5284 12955 5287
rect 13262 5284 13268 5296
rect 12943 5256 13268 5284
rect 12943 5253 12955 5256
rect 12897 5247 12955 5253
rect 13262 5244 13268 5256
rect 13320 5244 13326 5296
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 10100 5188 11897 5216
rect 10100 5176 10106 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12023 5188 13185 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 13173 5185 13185 5188
rect 13219 5216 13231 5219
rect 13446 5216 13452 5228
rect 13219 5188 13452 5216
rect 13219 5185 13231 5188
rect 13173 5179 13231 5185
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 6328 5120 6684 5148
rect 6328 5108 6334 5120
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 8202 5148 8208 5160
rect 7340 5120 8208 5148
rect 7340 5108 7346 5120
rect 8202 5108 8208 5120
rect 8260 5148 8266 5160
rect 10318 5148 10324 5160
rect 8260 5120 10324 5148
rect 8260 5108 8266 5120
rect 10318 5108 10324 5120
rect 10376 5148 10382 5160
rect 11701 5151 11759 5157
rect 11701 5148 11713 5151
rect 10376 5120 11713 5148
rect 10376 5108 10382 5120
rect 11701 5117 11713 5120
rect 11747 5117 11759 5151
rect 11701 5111 11759 5117
rect 11793 5151 11851 5157
rect 11793 5117 11805 5151
rect 11839 5117 11851 5151
rect 11793 5111 11851 5117
rect 8478 5080 8484 5092
rect 5920 5052 8484 5080
rect 8478 5040 8484 5052
rect 8536 5040 8542 5092
rect 10226 5040 10232 5092
rect 10284 5080 10290 5092
rect 11808 5080 11836 5111
rect 10284 5052 11836 5080
rect 10284 5040 10290 5052
rect 5169 5015 5227 5021
rect 5169 4981 5181 5015
rect 5215 4981 5227 5015
rect 5169 4975 5227 4981
rect 13354 4972 13360 5024
rect 13412 4972 13418 5024
rect 1104 4922 13800 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 13800 4922
rect 1104 4848 13800 4870
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 3418 4808 3424 4820
rect 2280 4780 3424 4808
rect 2280 4768 2286 4780
rect 3418 4768 3424 4780
rect 3476 4808 3482 4820
rect 5718 4808 5724 4820
rect 3476 4780 5724 4808
rect 3476 4768 3482 4780
rect 5718 4768 5724 4780
rect 5776 4768 5782 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 5902 4808 5908 4820
rect 5859 4780 5908 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 6086 4768 6092 4820
rect 6144 4768 6150 4820
rect 9490 4768 9496 4820
rect 9548 4768 9554 4820
rect 10597 4811 10655 4817
rect 10597 4777 10609 4811
rect 10643 4808 10655 4811
rect 10870 4808 10876 4820
rect 10643 4780 10876 4808
rect 10643 4777 10655 4780
rect 10597 4771 10655 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 5534 4700 5540 4752
rect 5592 4740 5598 4752
rect 6733 4743 6791 4749
rect 6733 4740 6745 4743
rect 5592 4712 6745 4740
rect 5592 4700 5598 4712
rect 6733 4709 6745 4712
rect 6779 4709 6791 4743
rect 6733 4703 6791 4709
rect 2958 4632 2964 4684
rect 3016 4632 3022 4684
rect 3142 4632 3148 4684
rect 3200 4632 3206 4684
rect 7834 4632 7840 4684
rect 7892 4672 7898 4684
rect 9217 4675 9275 4681
rect 9217 4672 9229 4675
rect 7892 4644 9229 4672
rect 7892 4632 7898 4644
rect 9217 4641 9229 4644
rect 9263 4641 9275 4675
rect 9217 4635 9275 4641
rect 842 4564 848 4616
rect 900 4604 906 4616
rect 1489 4607 1547 4613
rect 1489 4604 1501 4607
rect 900 4576 1501 4604
rect 900 4564 906 4576
rect 1489 4573 1501 4576
rect 1535 4573 1547 4607
rect 1489 4567 1547 4573
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4604 2099 4607
rect 2498 4604 2504 4616
rect 2087 4576 2504 4604
rect 2087 4573 2099 4576
rect 2041 4567 2099 4573
rect 2498 4564 2504 4576
rect 2556 4604 2562 4616
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2556 4576 2881 4604
rect 2556 4564 2562 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 4982 4564 4988 4616
rect 5040 4604 5046 4616
rect 5721 4607 5779 4613
rect 5721 4604 5733 4607
rect 5040 4576 5733 4604
rect 5040 4564 5046 4576
rect 5721 4573 5733 4576
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 5905 4607 5963 4613
rect 5905 4573 5917 4607
rect 5951 4604 5963 4607
rect 5994 4604 6000 4616
rect 5951 4576 6000 4604
rect 5951 4573 5963 4576
rect 5905 4567 5963 4573
rect 5994 4564 6000 4576
rect 6052 4564 6058 4616
rect 6362 4564 6368 4616
rect 6420 4604 6426 4616
rect 6549 4607 6607 4613
rect 6549 4604 6561 4607
rect 6420 4576 6561 4604
rect 6420 4564 6426 4576
rect 6549 4573 6561 4576
rect 6595 4604 6607 4607
rect 8846 4604 8852 4616
rect 6595 4576 8852 4604
rect 6595 4573 6607 4576
rect 6549 4567 6607 4573
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4573 9183 4607
rect 9232 4604 9260 4635
rect 10226 4604 10232 4616
rect 9232 4576 10232 4604
rect 9125 4567 9183 4573
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 5810 4536 5816 4548
rect 5408 4508 5816 4536
rect 5408 4496 5414 4508
rect 5810 4496 5816 4508
rect 5868 4536 5874 4548
rect 6273 4539 6331 4545
rect 6273 4536 6285 4539
rect 5868 4508 6285 4536
rect 5868 4496 5874 4508
rect 6273 4505 6285 4508
rect 6319 4505 6331 4539
rect 6273 4499 6331 4505
rect 6457 4539 6515 4545
rect 6457 4505 6469 4539
rect 6503 4536 6515 4539
rect 6638 4536 6644 4548
rect 6503 4508 6644 4536
rect 6503 4505 6515 4508
rect 6457 4499 6515 4505
rect 6638 4496 6644 4508
rect 6696 4536 6702 4548
rect 7006 4536 7012 4548
rect 6696 4508 7012 4536
rect 6696 4496 6702 4508
rect 7006 4496 7012 4508
rect 7064 4496 7070 4548
rect 8294 4496 8300 4548
rect 8352 4536 8358 4548
rect 9140 4536 9168 4567
rect 10226 4564 10232 4576
rect 10284 4564 10290 4616
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 8352 4508 9168 4536
rect 8352 4496 8358 4508
rect 9214 4496 9220 4548
rect 9272 4536 9278 4548
rect 10413 4539 10471 4545
rect 10413 4536 10425 4539
rect 9272 4508 10425 4536
rect 9272 4496 9278 4508
rect 10413 4505 10425 4508
rect 10459 4505 10471 4539
rect 10413 4499 10471 4505
rect 2498 4428 2504 4480
rect 2556 4428 2562 4480
rect 13262 4428 13268 4480
rect 13320 4428 13326 4480
rect 1104 4378 13800 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 13800 4378
rect 1104 4304 13800 4326
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 9033 4267 9091 4273
rect 9033 4264 9045 4267
rect 8352 4236 9045 4264
rect 8352 4224 8358 4236
rect 9033 4233 9045 4236
rect 9079 4264 9091 4267
rect 9858 4264 9864 4276
rect 9079 4236 9864 4264
rect 9079 4233 9091 4236
rect 9033 4227 9091 4233
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 10042 4224 10048 4276
rect 10100 4224 10106 4276
rect 2498 4156 2504 4208
rect 2556 4196 2562 4208
rect 2593 4199 2651 4205
rect 2593 4196 2605 4199
rect 2556 4168 2605 4196
rect 2556 4156 2562 4168
rect 2593 4165 2605 4168
rect 2639 4165 2651 4199
rect 3970 4196 3976 4208
rect 3818 4168 3976 4196
rect 2593 4159 2651 4165
rect 3970 4156 3976 4168
rect 4028 4156 4034 4208
rect 4341 4199 4399 4205
rect 4341 4165 4353 4199
rect 4387 4196 4399 4199
rect 5442 4196 5448 4208
rect 4387 4168 5448 4196
rect 4387 4165 4399 4168
rect 4341 4159 4399 4165
rect 5442 4156 5448 4168
rect 5500 4156 5506 4208
rect 7101 4199 7159 4205
rect 7101 4196 7113 4199
rect 6932 4168 7113 4196
rect 5810 4088 5816 4140
rect 5868 4088 5874 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 6932 4128 6960 4168
rect 7101 4165 7113 4168
rect 7147 4196 7159 4199
rect 7834 4196 7840 4208
rect 7147 4168 7840 4196
rect 7147 4165 7159 4168
rect 7101 4159 7159 4165
rect 7834 4156 7840 4168
rect 7892 4156 7898 4208
rect 10060 4196 10088 4224
rect 8956 4168 9168 4196
rect 6595 4100 6960 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 7006 4088 7012 4140
rect 7064 4088 7070 4140
rect 7282 4088 7288 4140
rect 7340 4088 7346 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7484 4100 7665 4128
rect 2314 4020 2320 4072
rect 2372 4020 2378 4072
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 5721 4063 5779 4069
rect 5721 4060 5733 4063
rect 5592 4032 5733 4060
rect 5592 4020 5598 4032
rect 5721 4029 5733 4032
rect 5767 4029 5779 4063
rect 5721 4023 5779 4029
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 6181 3995 6239 4001
rect 6181 3961 6193 3995
rect 6227 3992 6239 3995
rect 6656 3992 6684 4023
rect 6914 4020 6920 4072
rect 6972 4020 6978 4072
rect 7024 4060 7052 4088
rect 7484 4060 7512 4100
rect 7653 4097 7665 4100
rect 7699 4128 7711 4131
rect 7742 4128 7748 4140
rect 7699 4100 7748 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 8573 4131 8631 4137
rect 8573 4097 8585 4131
rect 8619 4128 8631 4131
rect 8956 4128 8984 4168
rect 8619 4100 8984 4128
rect 9140 4128 9168 4168
rect 9876 4168 10088 4196
rect 10137 4199 10195 4205
rect 9876 4128 9904 4168
rect 10137 4165 10149 4199
rect 10183 4196 10195 4199
rect 10870 4196 10876 4208
rect 10183 4168 10876 4196
rect 10183 4165 10195 4168
rect 10137 4159 10195 4165
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 9140 4100 9904 4128
rect 8619 4097 8631 4100
rect 8573 4091 8631 4097
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 10255 4131 10313 4137
rect 10255 4128 10267 4131
rect 10045 4091 10103 4097
rect 10152 4100 10267 4128
rect 7024 4032 7512 4060
rect 7561 4063 7619 4069
rect 7561 4029 7573 4063
rect 7607 4029 7619 4063
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 7561 4023 7619 4029
rect 7668 4032 9137 4060
rect 7576 3992 7604 4023
rect 6227 3964 7604 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 6546 3884 6552 3936
rect 6604 3924 6610 3936
rect 7009 3927 7067 3933
rect 7009 3924 7021 3927
rect 6604 3896 7021 3924
rect 6604 3884 6610 3896
rect 7009 3893 7021 3896
rect 7055 3893 7067 3927
rect 7009 3887 7067 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7668 3924 7696 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 8021 3995 8079 4001
rect 8021 3961 8033 3995
rect 8067 3992 8079 3995
rect 9030 3992 9036 4004
rect 8067 3964 9036 3992
rect 8067 3961 8079 3964
rect 8021 3955 8079 3961
rect 9030 3952 9036 3964
rect 9088 3952 9094 4004
rect 9140 3992 9168 4023
rect 9214 4020 9220 4072
rect 9272 4020 9278 4072
rect 9858 4020 9864 4072
rect 9916 4060 9922 4072
rect 10060 4060 10088 4091
rect 9916 4032 10088 4060
rect 9916 4020 9922 4032
rect 10152 3992 10180 4100
rect 10255 4097 10267 4100
rect 10301 4128 10313 4131
rect 10778 4128 10784 4140
rect 10301 4100 10784 4128
rect 10301 4097 10313 4100
rect 10255 4091 10313 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10244 4032 10425 4060
rect 10244 4004 10272 4032
rect 10413 4029 10425 4032
rect 10459 4029 10471 4063
rect 10413 4023 10471 4029
rect 9140 3964 10180 3992
rect 10226 3952 10232 4004
rect 10284 3952 10290 4004
rect 7156 3896 7696 3924
rect 7156 3884 7162 3896
rect 7742 3884 7748 3936
rect 7800 3924 7806 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 7800 3896 8401 3924
rect 7800 3884 7806 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 8570 3884 8576 3936
rect 8628 3924 8634 3936
rect 8665 3927 8723 3933
rect 8665 3924 8677 3927
rect 8628 3896 8677 3924
rect 8628 3884 8634 3896
rect 8665 3893 8677 3896
rect 8711 3893 8723 3927
rect 8665 3887 8723 3893
rect 9582 3884 9588 3936
rect 9640 3924 9646 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9640 3896 9781 3924
rect 9640 3884 9646 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 9769 3887 9827 3893
rect 1104 3834 13800 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 13800 3834
rect 1104 3760 13800 3782
rect 2406 3720 2412 3732
rect 1412 3692 2412 3720
rect 1412 3593 1440 3692
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 1397 3587 1455 3593
rect 1397 3553 1409 3587
rect 1443 3553 1455 3587
rect 1397 3547 1455 3553
rect 1670 3544 1676 3596
rect 1728 3544 1734 3596
rect 2406 3544 2412 3596
rect 2464 3584 2470 3596
rect 5261 3587 5319 3593
rect 5261 3584 5273 3587
rect 2464 3556 5273 3584
rect 2464 3544 2470 3556
rect 5261 3553 5273 3556
rect 5307 3553 5319 3587
rect 5261 3547 5319 3553
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 7340 3556 7604 3584
rect 7340 3544 7346 3556
rect 3418 3476 3424 3528
rect 3476 3476 3482 3528
rect 7576 3525 7604 3556
rect 9306 3544 9312 3596
rect 9364 3544 9370 3596
rect 9582 3544 9588 3596
rect 9640 3544 9646 3596
rect 10226 3544 10232 3596
rect 10284 3584 10290 3596
rect 11333 3587 11391 3593
rect 11333 3584 11345 3587
rect 10284 3556 11345 3584
rect 10284 3544 10290 3556
rect 11333 3553 11345 3556
rect 11379 3553 11391 3587
rect 11333 3547 11391 3553
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 7742 3476 7748 3528
rect 7800 3476 7806 3528
rect 7834 3476 7840 3528
rect 7892 3476 7898 3528
rect 3970 3448 3976 3460
rect 2898 3420 3976 3448
rect 3970 3408 3976 3420
rect 4028 3408 4034 3460
rect 5534 3408 5540 3460
rect 5592 3408 5598 3460
rect 7190 3448 7196 3460
rect 6762 3420 7196 3448
rect 7190 3408 7196 3420
rect 7248 3408 7254 3460
rect 10594 3408 10600 3460
rect 10652 3408 10658 3460
rect 7374 3340 7380 3392
rect 7432 3340 7438 3392
rect 1104 3290 13800 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 13800 3290
rect 1104 3216 13800 3238
rect 5534 3136 5540 3188
rect 5592 3176 5598 3188
rect 6365 3179 6423 3185
rect 6365 3176 6377 3179
rect 5592 3148 6377 3176
rect 5592 3136 5598 3148
rect 6365 3145 6377 3148
rect 6411 3145 6423 3179
rect 7190 3176 7196 3188
rect 6365 3139 6423 3145
rect 6472 3148 7196 3176
rect 2590 3068 2596 3120
rect 2648 3108 2654 3120
rect 2685 3111 2743 3117
rect 2685 3108 2697 3111
rect 2648 3080 2697 3108
rect 2648 3068 2654 3080
rect 2685 3077 2697 3080
rect 2731 3077 2743 3111
rect 3970 3108 3976 3120
rect 3910 3080 3976 3108
rect 2685 3071 2743 3077
rect 3970 3068 3976 3080
rect 4028 3108 4034 3120
rect 6472 3108 6500 3148
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 7484 3148 9904 3176
rect 4028 3080 6500 3108
rect 6641 3111 6699 3117
rect 4028 3068 4034 3080
rect 6641 3077 6653 3111
rect 6687 3108 6699 3111
rect 7374 3108 7380 3120
rect 6687 3080 7380 3108
rect 6687 3077 6699 3080
rect 6641 3071 6699 3077
rect 7374 3068 7380 3080
rect 7432 3068 7438 3120
rect 7484 3117 7512 3148
rect 7469 3111 7527 3117
rect 7469 3077 7481 3111
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 8570 3068 8576 3120
rect 8628 3068 8634 3120
rect 9876 3108 9904 3148
rect 9950 3136 9956 3188
rect 10008 3176 10014 3188
rect 10229 3179 10287 3185
rect 10229 3176 10241 3179
rect 10008 3148 10241 3176
rect 10008 3136 10014 3148
rect 10229 3145 10241 3148
rect 10275 3145 10287 3179
rect 10229 3139 10287 3145
rect 10594 3136 10600 3188
rect 10652 3136 10658 3188
rect 10612 3108 10640 3136
rect 9798 3080 10640 3108
rect 10873 3111 10931 3117
rect 10873 3077 10885 3111
rect 10919 3108 10931 3111
rect 13262 3108 13268 3120
rect 10919 3080 13268 3108
rect 10919 3077 10931 3080
rect 10873 3071 10931 3077
rect 13262 3068 13268 3080
rect 13320 3068 13326 3120
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 6546 3000 6552 3052
rect 6604 3000 6610 3052
rect 6914 3049 6920 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 6733 3003 6791 3009
rect 6871 3043 6920 3049
rect 6871 3009 6883 3043
rect 6917 3009 6920 3043
rect 6871 3003 6920 3009
rect 4157 2975 4215 2981
rect 4157 2941 4169 2975
rect 4203 2972 4215 2975
rect 6362 2972 6368 2984
rect 4203 2944 6368 2972
rect 4203 2941 4215 2944
rect 4157 2935 4215 2941
rect 6362 2932 6368 2944
rect 6420 2932 6426 2984
rect 6748 2972 6776 3003
rect 6914 3000 6920 3003
rect 6972 3000 6978 3052
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7282 3040 7288 3052
rect 7055 3012 7288 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 10229 3043 10287 3049
rect 10229 3040 10241 3043
rect 10152 3012 10241 3040
rect 10152 2984 10180 3012
rect 10229 3009 10241 3012
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10376 3012 10425 3040
rect 10376 3000 10382 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 8202 2972 8208 2984
rect 6748 2944 8208 2972
rect 8202 2932 8208 2944
rect 8260 2932 8266 2984
rect 8297 2975 8355 2981
rect 8297 2941 8309 2975
rect 8343 2972 8355 2975
rect 9306 2972 9312 2984
rect 8343 2944 9312 2972
rect 8343 2941 8355 2944
rect 8297 2935 8355 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 10045 2975 10103 2981
rect 10045 2941 10057 2975
rect 10091 2972 10103 2975
rect 10134 2972 10140 2984
rect 10091 2944 10140 2972
rect 10091 2941 10103 2944
rect 10045 2935 10103 2941
rect 10134 2932 10140 2944
rect 10192 2932 10198 2984
rect 1104 2746 13800 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 13800 2746
rect 1104 2672 13800 2694
rect 7190 2456 7196 2508
rect 7248 2496 7254 2508
rect 7248 2468 8800 2496
rect 7248 2456 7254 2468
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7742 2428 7748 2440
rect 7515 2400 7748 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8772 2437 8800 2468
rect 8113 2431 8171 2437
rect 8113 2428 8125 2431
rect 7892 2400 8125 2428
rect 7892 2388 7898 2400
rect 8113 2397 8125 2400
rect 8159 2397 8171 2431
rect 8113 2391 8171 2397
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 8757 2391 8815 2397
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7285 2295 7343 2301
rect 7285 2292 7297 2295
rect 7156 2264 7297 2292
rect 7156 2252 7162 2264
rect 7285 2261 7297 2264
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 7742 2252 7748 2304
rect 7800 2292 7806 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7800 2264 7941 2292
rect 7800 2252 7806 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 8386 2252 8392 2304
rect 8444 2292 8450 2304
rect 8573 2295 8631 2301
rect 8573 2292 8585 2295
rect 8444 2264 8585 2292
rect 8444 2252 8450 2264
rect 8573 2261 8585 2264
rect 8619 2261 8631 2295
rect 8573 2255 8631 2261
rect 1104 2202 13800 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 13800 2202
rect 1104 2128 13800 2150
<< via1 >>
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 9680 14560 9732 14612
rect 5816 14424 5868 14476
rect 6368 14356 6420 14408
rect 6092 14288 6144 14340
rect 7104 14356 7156 14408
rect 8392 14356 8444 14408
rect 10324 14356 10376 14408
rect 5816 14220 5868 14272
rect 6828 14220 6880 14272
rect 7840 14220 7892 14272
rect 8668 14263 8720 14272
rect 8668 14229 8677 14263
rect 8677 14229 8711 14263
rect 8711 14229 8720 14263
rect 8668 14220 8720 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 8024 14016 8076 14068
rect 7840 13948 7892 14000
rect 5448 13855 5500 13864
rect 5448 13821 5457 13855
rect 5457 13821 5491 13855
rect 5491 13821 5500 13855
rect 5448 13812 5500 13821
rect 5540 13744 5592 13796
rect 5908 13719 5960 13728
rect 5908 13685 5917 13719
rect 5917 13685 5951 13719
rect 5951 13685 5960 13719
rect 5908 13676 5960 13685
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7012 13880 7064 13889
rect 9404 13880 9456 13932
rect 9772 13880 9824 13932
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 10692 13880 10744 13932
rect 6828 13855 6880 13864
rect 6828 13821 6837 13855
rect 6837 13821 6871 13855
rect 6871 13821 6880 13855
rect 6828 13812 6880 13821
rect 8484 13744 8536 13796
rect 9956 13855 10008 13864
rect 9956 13821 9965 13855
rect 9965 13821 9999 13855
rect 9999 13821 10008 13855
rect 9956 13812 10008 13821
rect 6920 13676 6972 13728
rect 7196 13719 7248 13728
rect 7196 13685 7205 13719
rect 7205 13685 7239 13719
rect 7239 13685 7248 13719
rect 7196 13676 7248 13685
rect 8760 13676 8812 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 5448 13472 5500 13524
rect 5908 13472 5960 13524
rect 7012 13472 7064 13524
rect 7288 13472 7340 13524
rect 4804 13404 4856 13456
rect 5632 13404 5684 13456
rect 848 13268 900 13320
rect 4620 13336 4672 13388
rect 5816 13336 5868 13388
rect 9404 13404 9456 13456
rect 5448 13268 5500 13320
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 5724 13311 5776 13320
rect 5724 13277 5733 13311
rect 5733 13277 5767 13311
rect 5767 13277 5776 13311
rect 5724 13268 5776 13277
rect 7840 13311 7892 13320
rect 7840 13277 7849 13311
rect 7849 13277 7883 13311
rect 7883 13277 7892 13311
rect 7840 13268 7892 13277
rect 10692 13379 10744 13388
rect 10692 13345 10701 13379
rect 10701 13345 10735 13379
rect 10735 13345 10744 13379
rect 10692 13336 10744 13345
rect 8668 13268 8720 13320
rect 5264 13200 5316 13252
rect 6368 13200 6420 13252
rect 7564 13200 7616 13252
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 3884 13175 3936 13184
rect 3884 13141 3893 13175
rect 3893 13141 3927 13175
rect 3927 13141 3936 13175
rect 3884 13132 3936 13141
rect 5448 13132 5500 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 8852 13132 8904 13184
rect 10508 13200 10560 13252
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 2688 12928 2740 12980
rect 5632 12928 5684 12980
rect 6092 12928 6144 12980
rect 3792 12860 3844 12912
rect 4896 12860 4948 12912
rect 5724 12860 5776 12912
rect 6644 12903 6696 12912
rect 6644 12869 6653 12903
rect 6653 12869 6687 12903
rect 6687 12869 6696 12903
rect 6644 12860 6696 12869
rect 8484 12971 8536 12980
rect 8484 12937 8493 12971
rect 8493 12937 8527 12971
rect 8527 12937 8536 12971
rect 8484 12928 8536 12937
rect 9772 12971 9824 12980
rect 9772 12937 9781 12971
rect 9781 12937 9815 12971
rect 9815 12937 9824 12971
rect 9772 12928 9824 12937
rect 8024 12903 8076 12912
rect 8024 12869 8033 12903
rect 8033 12869 8067 12903
rect 8067 12869 8076 12903
rect 8024 12860 8076 12869
rect 8668 12860 8720 12912
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5356 12792 5408 12844
rect 5448 12792 5500 12844
rect 2872 12767 2924 12776
rect 2872 12733 2881 12767
rect 2881 12733 2915 12767
rect 2915 12733 2924 12767
rect 2872 12724 2924 12733
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 4712 12724 4764 12776
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 5816 12767 5868 12776
rect 5816 12733 5825 12767
rect 5825 12733 5859 12767
rect 5859 12733 5868 12767
rect 5816 12724 5868 12733
rect 6368 12792 6420 12844
rect 7012 12792 7064 12844
rect 7932 12792 7984 12844
rect 8852 12792 8904 12844
rect 10232 12792 10284 12844
rect 10508 12860 10560 12912
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 10048 12767 10100 12776
rect 10048 12733 10057 12767
rect 10057 12733 10091 12767
rect 10091 12733 10100 12767
rect 10048 12724 10100 12733
rect 6460 12656 6512 12708
rect 6920 12656 6972 12708
rect 9956 12656 10008 12708
rect 4620 12588 4672 12640
rect 7104 12588 7156 12640
rect 9404 12588 9456 12640
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 3700 12384 3752 12436
rect 4896 12384 4948 12436
rect 5356 12384 5408 12436
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 2688 12248 2740 12300
rect 1768 12223 1820 12232
rect 1768 12189 1777 12223
rect 1777 12189 1811 12223
rect 1811 12189 1820 12223
rect 1768 12180 1820 12189
rect 4160 12316 4212 12368
rect 4988 12316 5040 12368
rect 7012 12384 7064 12436
rect 10048 12384 10100 12436
rect 2872 12248 2924 12300
rect 3976 12248 4028 12300
rect 2964 12112 3016 12164
rect 3516 12223 3568 12232
rect 3516 12189 3525 12223
rect 3525 12189 3559 12223
rect 3559 12189 3568 12223
rect 3516 12180 3568 12189
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 5908 12248 5960 12300
rect 6920 12248 6972 12300
rect 7288 12359 7340 12368
rect 7288 12325 7297 12359
rect 7297 12325 7331 12359
rect 7331 12325 7340 12359
rect 7288 12316 7340 12325
rect 11796 12316 11848 12368
rect 8024 12180 8076 12232
rect 9588 12248 9640 12300
rect 10876 12248 10928 12300
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 10232 12223 10284 12232
rect 10232 12189 10241 12223
rect 10241 12189 10275 12223
rect 10275 12189 10284 12223
rect 10232 12180 10284 12189
rect 2596 12044 2648 12096
rect 3700 12112 3752 12164
rect 4804 12112 4856 12164
rect 6000 12112 6052 12164
rect 7564 12155 7616 12164
rect 7564 12121 7573 12155
rect 7573 12121 7607 12155
rect 7607 12121 7616 12155
rect 7564 12112 7616 12121
rect 7932 12112 7984 12164
rect 6552 12044 6604 12096
rect 7104 12044 7156 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 1400 11840 1452 11892
rect 1768 11840 1820 11892
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 6920 11840 6972 11892
rect 7196 11840 7248 11892
rect 9220 11840 9272 11892
rect 9496 11840 9548 11892
rect 1584 11772 1636 11824
rect 940 11636 992 11688
rect 1952 11543 2004 11552
rect 1952 11509 1961 11543
rect 1961 11509 1995 11543
rect 1995 11509 2004 11543
rect 1952 11500 2004 11509
rect 2688 11772 2740 11824
rect 4804 11772 4856 11824
rect 7472 11772 7524 11824
rect 2504 11747 2556 11756
rect 2504 11713 2513 11747
rect 2513 11713 2547 11747
rect 2547 11713 2556 11747
rect 2504 11704 2556 11713
rect 4896 11704 4948 11756
rect 5448 11704 5500 11756
rect 2964 11636 3016 11688
rect 4712 11636 4764 11688
rect 5356 11636 5408 11688
rect 5724 11747 5776 11756
rect 5724 11713 5733 11747
rect 5733 11713 5767 11747
rect 5767 11713 5776 11747
rect 5724 11704 5776 11713
rect 6920 11704 6972 11756
rect 7564 11704 7616 11756
rect 7840 11747 7892 11756
rect 7840 11713 7849 11747
rect 7849 11713 7883 11747
rect 7883 11713 7892 11747
rect 7840 11704 7892 11713
rect 9404 11772 9456 11824
rect 10416 11704 10468 11756
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 7104 11636 7156 11688
rect 9312 11679 9364 11688
rect 9312 11645 9321 11679
rect 9321 11645 9355 11679
rect 9355 11645 9364 11679
rect 9312 11636 9364 11645
rect 6460 11611 6512 11620
rect 6460 11577 6469 11611
rect 6469 11577 6503 11611
rect 6503 11577 6512 11611
rect 6460 11568 6512 11577
rect 4712 11500 4764 11552
rect 5540 11500 5592 11552
rect 7564 11500 7616 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 3240 11296 3292 11348
rect 4712 11296 4764 11348
rect 3516 11228 3568 11280
rect 3976 11228 4028 11280
rect 9312 11296 9364 11348
rect 11152 11228 11204 11280
rect 3240 11160 3292 11212
rect 5540 11203 5592 11212
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 1952 11092 2004 11144
rect 2504 11135 2556 11144
rect 2504 11101 2513 11135
rect 2513 11101 2547 11135
rect 2547 11101 2556 11135
rect 2504 11092 2556 11101
rect 4068 11092 4120 11144
rect 4712 11092 4764 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 9036 11203 9088 11212
rect 9036 11169 9045 11203
rect 9045 11169 9079 11203
rect 9079 11169 9088 11203
rect 9036 11160 9088 11169
rect 8024 11092 8076 11144
rect 9496 11092 9548 11144
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 4620 11024 4672 11076
rect 5540 11024 5592 11076
rect 6000 11024 6052 11076
rect 7840 11024 7892 11076
rect 11704 11067 11756 11076
rect 11704 11033 11713 11067
rect 11713 11033 11747 11067
rect 11747 11033 11756 11067
rect 11704 11024 11756 11033
rect 12716 11024 12768 11076
rect 13176 11024 13228 11076
rect 11888 10956 11940 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3884 10752 3936 10804
rect 4620 10752 4672 10804
rect 5724 10795 5776 10804
rect 5724 10761 5733 10795
rect 5733 10761 5767 10795
rect 5767 10761 5776 10795
rect 5724 10752 5776 10761
rect 7104 10752 7156 10804
rect 11704 10752 11756 10804
rect 6368 10684 6420 10736
rect 7564 10659 7616 10668
rect 7564 10625 7573 10659
rect 7573 10625 7607 10659
rect 7607 10625 7616 10659
rect 7564 10616 7616 10625
rect 9128 10659 9180 10668
rect 9128 10625 9137 10659
rect 9137 10625 9171 10659
rect 9171 10625 9180 10659
rect 9128 10616 9180 10625
rect 9588 10616 9640 10668
rect 11152 10659 11204 10668
rect 11152 10625 11161 10659
rect 11161 10625 11195 10659
rect 11195 10625 11204 10659
rect 11152 10616 11204 10625
rect 13176 10684 13228 10736
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 8576 10548 8628 10600
rect 11888 10616 11940 10668
rect 12256 10616 12308 10668
rect 11796 10591 11848 10600
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 12440 10548 12492 10600
rect 11888 10480 11940 10532
rect 9956 10412 10008 10464
rect 11428 10412 11480 10464
rect 12348 10412 12400 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 9036 10208 9088 10260
rect 1400 10072 1452 10124
rect 3700 10004 3752 10056
rect 8300 10047 8352 10056
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9220 10047 9272 10056
rect 9220 10013 9229 10047
rect 9229 10013 9263 10047
rect 9263 10013 9272 10047
rect 9220 10004 9272 10013
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 9496 9979 9548 9988
rect 9496 9945 9505 9979
rect 9505 9945 9539 9979
rect 9539 9945 9548 9979
rect 9496 9936 9548 9945
rect 11704 9979 11756 9988
rect 11704 9945 11713 9979
rect 11713 9945 11747 9979
rect 11747 9945 11756 9979
rect 11704 9936 11756 9945
rect 12716 9936 12768 9988
rect 13084 9936 13136 9988
rect 3700 9868 3752 9920
rect 8392 9911 8444 9920
rect 8392 9877 8401 9911
rect 8401 9877 8435 9911
rect 8435 9877 8444 9911
rect 8392 9868 8444 9877
rect 8760 9911 8812 9920
rect 8760 9877 8769 9911
rect 8769 9877 8803 9911
rect 8803 9877 8812 9911
rect 8760 9868 8812 9877
rect 9036 9868 9088 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 10324 9868 10376 9920
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 8760 9664 8812 9716
rect 9312 9664 9364 9716
rect 9496 9707 9548 9716
rect 9496 9673 9505 9707
rect 9505 9673 9539 9707
rect 9539 9673 9548 9707
rect 9496 9664 9548 9673
rect 11704 9664 11756 9716
rect 3976 9596 4028 9648
rect 6552 9596 6604 9648
rect 8576 9596 8628 9648
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 6092 9571 6144 9580
rect 6092 9537 6101 9571
rect 6101 9537 6135 9571
rect 6135 9537 6144 9571
rect 6092 9528 6144 9537
rect 6276 9528 6328 9580
rect 6460 9528 6512 9580
rect 1676 9503 1728 9512
rect 1676 9469 1685 9503
rect 1685 9469 1719 9503
rect 1719 9469 1728 9503
rect 1676 9460 1728 9469
rect 2228 9460 2280 9512
rect 3516 9503 3568 9512
rect 3516 9469 3525 9503
rect 3525 9469 3559 9503
rect 3559 9469 3568 9503
rect 3516 9460 3568 9469
rect 3976 9460 4028 9512
rect 5540 9460 5592 9512
rect 5816 9460 5868 9512
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 7012 9571 7064 9580
rect 7012 9537 7021 9571
rect 7021 9537 7055 9571
rect 7055 9537 7064 9571
rect 7012 9528 7064 9537
rect 7932 9528 7984 9580
rect 9588 9596 9640 9648
rect 9956 9639 10008 9648
rect 9956 9605 9965 9639
rect 9965 9605 9999 9639
rect 9999 9605 10008 9639
rect 9956 9596 10008 9605
rect 10876 9639 10928 9648
rect 10876 9605 10885 9639
rect 10885 9605 10919 9639
rect 10919 9605 10928 9639
rect 10876 9596 10928 9605
rect 12164 9664 12216 9716
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 8760 9503 8812 9512
rect 8760 9469 8769 9503
rect 8769 9469 8803 9503
rect 8803 9469 8812 9503
rect 8760 9460 8812 9469
rect 9864 9460 9916 9512
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 10324 9571 10376 9580
rect 10324 9537 10333 9571
rect 10333 9537 10367 9571
rect 10367 9537 10376 9571
rect 10324 9528 10376 9537
rect 10600 9571 10652 9580
rect 10600 9537 10609 9571
rect 10609 9537 10643 9571
rect 10643 9537 10652 9571
rect 10600 9528 10652 9537
rect 10692 9571 10744 9580
rect 10692 9537 10701 9571
rect 10701 9537 10735 9571
rect 10735 9537 10744 9571
rect 10692 9528 10744 9537
rect 2228 9324 2280 9376
rect 4804 9324 4856 9376
rect 5540 9324 5592 9376
rect 5908 9324 5960 9376
rect 8116 9324 8168 9376
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 13084 9596 13136 9648
rect 12624 9528 12676 9537
rect 13176 9571 13228 9580
rect 13176 9537 13185 9571
rect 13185 9537 13219 9571
rect 13219 9537 13228 9571
rect 13176 9528 13228 9537
rect 12164 9503 12216 9512
rect 12164 9469 12173 9503
rect 12173 9469 12207 9503
rect 12207 9469 12216 9503
rect 12164 9460 12216 9469
rect 13360 9435 13412 9444
rect 13360 9401 13369 9435
rect 13369 9401 13403 9435
rect 13403 9401 13412 9435
rect 13360 9392 13412 9401
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 1860 9120 1912 9172
rect 3516 9120 3568 9172
rect 2320 9052 2372 9104
rect 848 8916 900 8968
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 2596 8984 2648 9036
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 4712 9052 4764 9104
rect 5632 9120 5684 9172
rect 6092 9120 6144 9172
rect 6460 9163 6512 9172
rect 6460 9129 6469 9163
rect 6469 9129 6503 9163
rect 6503 9129 6512 9163
rect 6460 9120 6512 9129
rect 6828 9120 6880 9172
rect 8760 9163 8812 9172
rect 8760 9129 8769 9163
rect 8769 9129 8803 9163
rect 8803 9129 8812 9163
rect 8760 9120 8812 9129
rect 10048 9120 10100 9172
rect 11244 9120 11296 9172
rect 12164 9120 12216 9172
rect 5816 9052 5868 9104
rect 6184 9052 6236 9104
rect 4344 9027 4396 9036
rect 4344 8993 4353 9027
rect 4353 8993 4387 9027
rect 4387 8993 4396 9027
rect 4344 8984 4396 8993
rect 5724 8984 5776 9036
rect 4620 8916 4672 8968
rect 4804 8916 4856 8968
rect 3700 8848 3752 8900
rect 2136 8780 2188 8832
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 2964 8823 3016 8832
rect 2964 8789 2973 8823
rect 2973 8789 3007 8823
rect 3007 8789 3016 8823
rect 2964 8780 3016 8789
rect 3056 8780 3108 8832
rect 4344 8848 4396 8900
rect 5356 8959 5408 8968
rect 5356 8925 5365 8959
rect 5365 8925 5399 8959
rect 5399 8925 5408 8959
rect 5356 8916 5408 8925
rect 5908 8916 5960 8968
rect 6276 8984 6328 9036
rect 6736 8984 6788 9036
rect 6368 8848 6420 8900
rect 6644 8916 6696 8968
rect 6736 8848 6788 8900
rect 8944 9052 8996 9104
rect 8392 8984 8444 9036
rect 8668 8984 8720 9036
rect 5356 8780 5408 8832
rect 5540 8780 5592 8832
rect 6276 8823 6328 8832
rect 6276 8789 6285 8823
rect 6285 8789 6319 8823
rect 6319 8789 6328 8823
rect 6276 8780 6328 8789
rect 6460 8780 6512 8832
rect 6828 8780 6880 8832
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 8760 8916 8812 8968
rect 8852 8916 8904 8968
rect 8208 8891 8260 8900
rect 8208 8857 8217 8891
rect 8217 8857 8251 8891
rect 8251 8857 8260 8891
rect 8208 8848 8260 8857
rect 8944 8891 8996 8900
rect 8944 8857 8953 8891
rect 8953 8857 8987 8891
rect 8987 8857 8996 8891
rect 8944 8848 8996 8857
rect 9128 8916 9180 8968
rect 9588 8984 9640 9036
rect 11152 8916 11204 8968
rect 12532 8959 12584 8968
rect 12532 8925 12541 8959
rect 12541 8925 12575 8959
rect 12575 8925 12584 8959
rect 12532 8916 12584 8925
rect 12624 8959 12676 8968
rect 12624 8925 12633 8959
rect 12633 8925 12667 8959
rect 12667 8925 12676 8959
rect 12624 8916 12676 8925
rect 13084 8916 13136 8968
rect 11980 8848 12032 8900
rect 8116 8780 8168 8832
rect 9404 8780 9456 8832
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 12440 8823 12492 8832
rect 12440 8789 12449 8823
rect 12449 8789 12483 8823
rect 12483 8789 12492 8823
rect 12440 8780 12492 8789
rect 13360 8823 13412 8832
rect 13360 8789 13369 8823
rect 13369 8789 13403 8823
rect 13403 8789 13412 8823
rect 13360 8780 13412 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 1676 8576 1728 8628
rect 2596 8576 2648 8628
rect 5632 8576 5684 8628
rect 6092 8576 6144 8628
rect 2412 8508 2464 8560
rect 6552 8576 6604 8628
rect 7012 8576 7064 8628
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1768 8440 1820 8492
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 6368 8551 6420 8560
rect 6368 8517 6377 8551
rect 6377 8517 6411 8551
rect 6411 8517 6420 8551
rect 6368 8508 6420 8517
rect 2780 8304 2832 8356
rect 3332 8415 3384 8424
rect 3332 8381 3341 8415
rect 3341 8381 3375 8415
rect 3375 8381 3384 8415
rect 3332 8372 3384 8381
rect 3700 8304 3752 8356
rect 5724 8440 5776 8492
rect 6460 8440 6512 8492
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 8300 8576 8352 8628
rect 8944 8576 8996 8628
rect 9128 8619 9180 8628
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 12624 8576 12676 8628
rect 8208 8508 8260 8560
rect 6644 8440 6696 8449
rect 8116 8440 8168 8492
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 11060 8508 11112 8560
rect 11888 8508 11940 8560
rect 12808 8508 12860 8560
rect 9404 8440 9456 8492
rect 5356 8372 5408 8424
rect 8208 8372 8260 8424
rect 4528 8304 4580 8356
rect 5816 8304 5868 8356
rect 6184 8304 6236 8356
rect 8576 8372 8628 8424
rect 9220 8372 9272 8424
rect 11244 8372 11296 8424
rect 11428 8372 11480 8424
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 11888 8372 11940 8424
rect 12532 8372 12584 8424
rect 4068 8279 4120 8288
rect 4068 8245 4077 8279
rect 4077 8245 4111 8279
rect 4111 8245 4120 8279
rect 4068 8236 4120 8245
rect 5080 8236 5132 8288
rect 5632 8236 5684 8288
rect 6736 8236 6788 8288
rect 8668 8279 8720 8288
rect 8668 8245 8677 8279
rect 8677 8245 8711 8279
rect 8711 8245 8720 8279
rect 8668 8236 8720 8245
rect 8760 8236 8812 8288
rect 11152 8279 11204 8288
rect 11152 8245 11161 8279
rect 11161 8245 11195 8279
rect 11195 8245 11204 8279
rect 11152 8236 11204 8245
rect 13268 8279 13320 8288
rect 13268 8245 13277 8279
rect 13277 8245 13311 8279
rect 13311 8245 13320 8279
rect 13268 8236 13320 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 5356 8032 5408 8084
rect 5724 8032 5776 8084
rect 11152 8075 11204 8084
rect 11152 8041 11161 8075
rect 11161 8041 11195 8075
rect 11195 8041 11204 8075
rect 11152 8032 11204 8041
rect 11796 8032 11848 8084
rect 13360 8075 13412 8084
rect 13360 8041 13369 8075
rect 13369 8041 13403 8075
rect 13403 8041 13412 8075
rect 13360 8032 13412 8041
rect 2044 7871 2096 7880
rect 2044 7837 2053 7871
rect 2053 7837 2087 7871
rect 2087 7837 2096 7871
rect 2044 7828 2096 7837
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 3332 7896 3384 7948
rect 3792 7939 3844 7948
rect 3792 7905 3801 7939
rect 3801 7905 3835 7939
rect 3835 7905 3844 7939
rect 3792 7896 3844 7905
rect 4436 7896 4488 7948
rect 4620 7896 4672 7948
rect 2596 7828 2648 7880
rect 6460 7964 6512 8016
rect 8852 7964 8904 8016
rect 5632 7896 5684 7948
rect 6092 7896 6144 7948
rect 11060 7896 11112 7948
rect 5448 7828 5500 7880
rect 5540 7871 5592 7880
rect 5540 7837 5549 7871
rect 5549 7837 5583 7871
rect 5583 7837 5592 7871
rect 5540 7828 5592 7837
rect 4068 7760 4120 7812
rect 4712 7760 4764 7812
rect 5356 7760 5408 7812
rect 6552 7828 6604 7880
rect 8576 7828 8628 7880
rect 9220 7871 9272 7880
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 9588 7828 9640 7880
rect 11244 7871 11296 7880
rect 11244 7837 11253 7871
rect 11253 7837 11287 7871
rect 11287 7837 11296 7871
rect 11244 7828 11296 7837
rect 1860 7692 1912 7744
rect 2688 7735 2740 7744
rect 2688 7701 2697 7735
rect 2697 7701 2731 7735
rect 2731 7701 2740 7735
rect 2688 7692 2740 7701
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3332 7692 3384 7701
rect 4896 7692 4948 7744
rect 6828 7760 6880 7812
rect 11152 7760 11204 7812
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 11980 7871 12032 7880
rect 11980 7837 11989 7871
rect 11989 7837 12023 7871
rect 12023 7837 12032 7871
rect 11980 7828 12032 7837
rect 12072 7871 12124 7880
rect 12072 7837 12081 7871
rect 12081 7837 12115 7871
rect 12115 7837 12124 7871
rect 12072 7828 12124 7837
rect 6368 7735 6420 7744
rect 6368 7701 6377 7735
rect 6377 7701 6411 7735
rect 6411 7701 6420 7735
rect 6368 7692 6420 7701
rect 9496 7692 9548 7744
rect 11060 7692 11112 7744
rect 12256 7828 12308 7880
rect 12440 7828 12492 7880
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 12348 7735 12400 7744
rect 12348 7701 12357 7735
rect 12357 7701 12391 7735
rect 12391 7701 12400 7735
rect 12348 7692 12400 7701
rect 12624 7760 12676 7812
rect 13268 7828 13320 7880
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2504 7488 2556 7540
rect 2596 7488 2648 7540
rect 6920 7531 6972 7540
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 8760 7488 8812 7540
rect 2044 7420 2096 7472
rect 3884 7420 3936 7472
rect 5264 7420 5316 7472
rect 6368 7463 6420 7472
rect 6368 7429 6377 7463
rect 6377 7429 6411 7463
rect 6411 7429 6420 7463
rect 6368 7420 6420 7429
rect 6828 7420 6880 7472
rect 9220 7531 9272 7540
rect 9220 7497 9229 7531
rect 9229 7497 9263 7531
rect 9263 7497 9272 7531
rect 9220 7488 9272 7497
rect 9312 7488 9364 7540
rect 10600 7488 10652 7540
rect 12808 7488 12860 7540
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 2596 7352 2648 7361
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 3608 7395 3660 7404
rect 3608 7361 3617 7395
rect 3617 7361 3651 7395
rect 3651 7361 3660 7395
rect 3608 7352 3660 7361
rect 3792 7395 3844 7404
rect 3792 7361 3798 7395
rect 3798 7361 3844 7395
rect 3792 7352 3844 7361
rect 4436 7352 4488 7404
rect 5448 7352 5500 7404
rect 2688 7284 2740 7336
rect 5356 7284 5408 7336
rect 6184 7352 6236 7404
rect 7104 7352 7156 7404
rect 8852 7284 8904 7336
rect 9128 7395 9180 7404
rect 9128 7361 9137 7395
rect 9137 7361 9171 7395
rect 9171 7361 9180 7395
rect 9128 7352 9180 7361
rect 9312 7395 9364 7404
rect 9312 7361 9321 7395
rect 9321 7361 9355 7395
rect 9355 7361 9364 7395
rect 9312 7352 9364 7361
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 12900 7420 12952 7472
rect 9772 7395 9824 7404
rect 9772 7361 9781 7395
rect 9781 7361 9815 7395
rect 9815 7361 9824 7395
rect 9772 7352 9824 7361
rect 9864 7352 9916 7404
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 11428 7284 11480 7336
rect 11888 7327 11940 7336
rect 11888 7293 11897 7327
rect 11897 7293 11931 7327
rect 11931 7293 11940 7327
rect 11888 7284 11940 7293
rect 2964 7216 3016 7268
rect 3240 7148 3292 7200
rect 9496 7191 9548 7200
rect 9496 7157 9505 7191
rect 9505 7157 9539 7191
rect 9539 7157 9548 7191
rect 9496 7148 9548 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3608 6944 3660 6996
rect 11888 6944 11940 6996
rect 2044 6851 2096 6860
rect 2044 6817 2053 6851
rect 2053 6817 2087 6851
rect 2087 6817 2096 6851
rect 2044 6808 2096 6817
rect 3148 6876 3200 6928
rect 3056 6851 3108 6860
rect 3056 6817 3065 6851
rect 3065 6817 3099 6851
rect 3099 6817 3108 6851
rect 3056 6808 3108 6817
rect 8852 6876 8904 6928
rect 10232 6876 10284 6928
rect 848 6740 900 6792
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 4344 6808 4396 6860
rect 8484 6851 8536 6860
rect 8484 6817 8493 6851
rect 8493 6817 8527 6851
rect 8527 6817 8536 6851
rect 8484 6808 8536 6817
rect 3792 6783 3844 6792
rect 3792 6749 3801 6783
rect 3801 6749 3835 6783
rect 3835 6749 3844 6783
rect 3792 6740 3844 6749
rect 3884 6783 3936 6792
rect 3884 6749 3894 6783
rect 3894 6749 3928 6783
rect 3928 6749 3936 6783
rect 3884 6740 3936 6749
rect 3148 6672 3200 6724
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 4160 6715 4212 6724
rect 4160 6681 4169 6715
rect 4169 6681 4203 6715
rect 4203 6681 4212 6715
rect 4160 6672 4212 6681
rect 3608 6604 3660 6656
rect 8208 6740 8260 6792
rect 9036 6808 9088 6860
rect 9772 6808 9824 6860
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 9680 6783 9732 6792
rect 9680 6749 9689 6783
rect 9689 6749 9723 6783
rect 9723 6749 9732 6783
rect 9680 6740 9732 6749
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 12348 6808 12400 6860
rect 12440 6851 12492 6860
rect 12440 6817 12449 6851
rect 12449 6817 12483 6851
rect 12483 6817 12492 6851
rect 12440 6808 12492 6817
rect 12624 6740 12676 6792
rect 9404 6647 9456 6656
rect 9404 6613 9413 6647
rect 9413 6613 9447 6647
rect 9447 6613 9456 6647
rect 9404 6604 9456 6613
rect 10416 6647 10468 6656
rect 10416 6613 10425 6647
rect 10425 6613 10459 6647
rect 10459 6613 10468 6647
rect 10416 6604 10468 6613
rect 12164 6715 12216 6724
rect 12164 6681 12173 6715
rect 12173 6681 12207 6715
rect 12207 6681 12216 6715
rect 12164 6672 12216 6681
rect 12256 6715 12308 6724
rect 12256 6681 12291 6715
rect 12291 6681 12308 6715
rect 12256 6672 12308 6681
rect 12440 6672 12492 6724
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 1676 6375 1728 6384
rect 1676 6341 1685 6375
rect 1685 6341 1719 6375
rect 1719 6341 1728 6375
rect 1676 6332 1728 6341
rect 2872 6400 2924 6452
rect 2504 6332 2556 6384
rect 940 6264 992 6316
rect 4344 6400 4396 6452
rect 4160 6332 4212 6384
rect 5356 6400 5408 6452
rect 6828 6400 6880 6452
rect 5448 6332 5500 6384
rect 4712 6264 4764 6316
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 2044 6239 2096 6248
rect 2044 6205 2053 6239
rect 2053 6205 2087 6239
rect 2087 6205 2096 6239
rect 2044 6196 2096 6205
rect 2412 6196 2464 6248
rect 3976 6196 4028 6248
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5816 6332 5868 6384
rect 8944 6443 8996 6452
rect 8944 6409 8953 6443
rect 8953 6409 8987 6443
rect 8987 6409 8996 6443
rect 8944 6400 8996 6409
rect 9404 6400 9456 6452
rect 10692 6400 10744 6452
rect 10784 6400 10836 6452
rect 12256 6400 12308 6452
rect 5356 6264 5408 6273
rect 5724 6264 5776 6316
rect 6460 6307 6512 6316
rect 6460 6273 6469 6307
rect 6469 6273 6503 6307
rect 6503 6273 6512 6307
rect 6460 6264 6512 6273
rect 5448 6196 5500 6248
rect 5540 6239 5592 6248
rect 5540 6205 5549 6239
rect 5549 6205 5583 6239
rect 5583 6205 5592 6239
rect 5540 6196 5592 6205
rect 6552 6196 6604 6248
rect 6736 6307 6788 6316
rect 6736 6273 6745 6307
rect 6745 6273 6779 6307
rect 6779 6273 6788 6307
rect 6736 6264 6788 6273
rect 6920 6264 6972 6316
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 7012 6196 7064 6248
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 2504 6060 2556 6112
rect 4804 6128 4856 6180
rect 8760 6375 8812 6384
rect 8760 6341 8769 6375
rect 8769 6341 8803 6375
rect 8803 6341 8812 6375
rect 8760 6332 8812 6341
rect 10416 6332 10468 6384
rect 11060 6375 11112 6384
rect 11060 6341 11069 6375
rect 11069 6341 11103 6375
rect 11103 6341 11112 6375
rect 11060 6332 11112 6341
rect 5540 6103 5592 6112
rect 5540 6069 5549 6103
rect 5549 6069 5583 6103
rect 5583 6069 5592 6103
rect 8116 6264 8168 6316
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 9036 6307 9088 6316
rect 9036 6273 9045 6307
rect 9045 6273 9079 6307
rect 9079 6273 9088 6307
rect 9036 6264 9088 6273
rect 8024 6171 8076 6180
rect 8024 6137 8033 6171
rect 8033 6137 8067 6171
rect 8067 6137 8076 6171
rect 8024 6128 8076 6137
rect 8944 6196 8996 6248
rect 10324 6264 10376 6316
rect 12440 6264 12492 6316
rect 9220 6196 9272 6248
rect 9496 6196 9548 6248
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 5540 6060 5592 6069
rect 9588 6128 9640 6180
rect 10140 6128 10192 6180
rect 9680 6060 9732 6112
rect 10692 6060 10744 6112
rect 11060 6060 11112 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3240 5899 3292 5908
rect 3240 5865 3249 5899
rect 3249 5865 3283 5899
rect 3283 5865 3292 5899
rect 3240 5856 3292 5865
rect 3608 5856 3660 5908
rect 3792 5788 3844 5840
rect 3056 5720 3108 5772
rect 848 5652 900 5704
rect 2136 5652 2188 5704
rect 2228 5652 2280 5704
rect 2044 5584 2096 5636
rect 2964 5584 3016 5636
rect 4804 5652 4856 5704
rect 5724 5788 5776 5840
rect 5908 5763 5960 5772
rect 5908 5729 5917 5763
rect 5917 5729 5951 5763
rect 5951 5729 5960 5763
rect 5908 5720 5960 5729
rect 6184 5831 6236 5840
rect 6184 5797 6193 5831
rect 6193 5797 6227 5831
rect 6227 5797 6236 5831
rect 6184 5788 6236 5797
rect 6736 5856 6788 5908
rect 8944 5856 8996 5908
rect 9312 5899 9364 5908
rect 9312 5865 9321 5899
rect 9321 5865 9355 5899
rect 9355 5865 9364 5899
rect 9312 5856 9364 5865
rect 12440 5856 12492 5908
rect 8208 5788 8260 5840
rect 8852 5788 8904 5840
rect 9128 5788 9180 5840
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 6644 5652 6696 5704
rect 6828 5652 6880 5704
rect 8024 5652 8076 5704
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8484 5720 8536 5772
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 8852 5652 8904 5704
rect 5448 5584 5500 5636
rect 9220 5584 9272 5636
rect 4804 5516 4856 5568
rect 5356 5516 5408 5568
rect 6552 5516 6604 5568
rect 8116 5516 8168 5568
rect 9404 5516 9456 5568
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 10692 5695 10744 5704
rect 10692 5661 10701 5695
rect 10701 5661 10735 5695
rect 10735 5661 10744 5695
rect 10692 5652 10744 5661
rect 11060 5695 11112 5704
rect 11060 5661 11069 5695
rect 11069 5661 11103 5695
rect 11103 5661 11112 5695
rect 11060 5652 11112 5661
rect 11152 5695 11204 5704
rect 11152 5661 11161 5695
rect 11161 5661 11195 5695
rect 11195 5661 11204 5695
rect 11152 5652 11204 5661
rect 12808 5652 12860 5704
rect 10048 5627 10100 5636
rect 10048 5593 10057 5627
rect 10057 5593 10091 5627
rect 10091 5593 10100 5627
rect 10048 5584 10100 5593
rect 9864 5516 9916 5568
rect 10232 5559 10284 5568
rect 10232 5525 10241 5559
rect 10241 5525 10275 5559
rect 10275 5525 10284 5559
rect 10232 5516 10284 5525
rect 10784 5584 10836 5636
rect 13452 5627 13504 5636
rect 13452 5593 13461 5627
rect 13461 5593 13495 5627
rect 13495 5593 13504 5627
rect 13452 5584 13504 5593
rect 12072 5516 12124 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2044 5312 2096 5364
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 848 5176 900 5228
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 11152 5312 11204 5364
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 6000 5244 6052 5296
rect 6460 5244 6512 5296
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 2228 5108 2280 5117
rect 3148 5151 3200 5160
rect 3148 5117 3157 5151
rect 3157 5117 3191 5151
rect 3191 5117 3200 5151
rect 3148 5108 3200 5117
rect 5448 5176 5500 5228
rect 5724 5176 5776 5228
rect 6092 5176 6144 5228
rect 6552 5219 6604 5228
rect 6552 5185 6561 5219
rect 6561 5185 6595 5219
rect 6595 5185 6604 5219
rect 6552 5176 6604 5185
rect 10692 5244 10744 5296
rect 5356 5108 5408 5160
rect 1676 4972 1728 5024
rect 2596 5015 2648 5024
rect 2596 4981 2605 5015
rect 2605 4981 2639 5015
rect 2639 4981 2648 5015
rect 2596 4972 2648 4981
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 5540 5040 5592 5092
rect 6276 5108 6328 5160
rect 10048 5176 10100 5228
rect 13268 5244 13320 5296
rect 13452 5176 13504 5228
rect 7288 5108 7340 5160
rect 8208 5108 8260 5160
rect 10324 5108 10376 5160
rect 8484 5040 8536 5092
rect 10232 5040 10284 5092
rect 13360 5015 13412 5024
rect 13360 4981 13369 5015
rect 13369 4981 13403 5015
rect 13403 4981 13412 5015
rect 13360 4972 13412 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2228 4768 2280 4820
rect 3424 4768 3476 4820
rect 5724 4768 5776 4820
rect 5908 4768 5960 4820
rect 6092 4811 6144 4820
rect 6092 4777 6101 4811
rect 6101 4777 6135 4811
rect 6135 4777 6144 4811
rect 6092 4768 6144 4777
rect 9496 4811 9548 4820
rect 9496 4777 9505 4811
rect 9505 4777 9539 4811
rect 9539 4777 9548 4811
rect 9496 4768 9548 4777
rect 10876 4768 10928 4820
rect 5540 4700 5592 4752
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 3148 4675 3200 4684
rect 3148 4641 3157 4675
rect 3157 4641 3191 4675
rect 3191 4641 3200 4675
rect 3148 4632 3200 4641
rect 7840 4632 7892 4684
rect 848 4564 900 4616
rect 2504 4564 2556 4616
rect 4988 4564 5040 4616
rect 6000 4564 6052 4616
rect 6368 4564 6420 4616
rect 8852 4564 8904 4616
rect 10232 4607 10284 4616
rect 5356 4496 5408 4548
rect 5816 4496 5868 4548
rect 6644 4496 6696 4548
rect 7012 4496 7064 4548
rect 8300 4496 8352 4548
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 9220 4496 9272 4548
rect 2504 4471 2556 4480
rect 2504 4437 2513 4471
rect 2513 4437 2547 4471
rect 2547 4437 2556 4471
rect 2504 4428 2556 4437
rect 13268 4471 13320 4480
rect 13268 4437 13277 4471
rect 13277 4437 13311 4471
rect 13311 4437 13320 4471
rect 13268 4428 13320 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 8300 4224 8352 4276
rect 9864 4224 9916 4276
rect 10048 4224 10100 4276
rect 2504 4156 2556 4208
rect 3976 4156 4028 4208
rect 5448 4156 5500 4208
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 7840 4156 7892 4208
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 2320 4063 2372 4072
rect 2320 4029 2329 4063
rect 2329 4029 2363 4063
rect 2363 4029 2372 4063
rect 2320 4020 2372 4029
rect 5540 4020 5592 4072
rect 6920 4063 6972 4072
rect 6920 4029 6929 4063
rect 6929 4029 6963 4063
rect 6963 4029 6972 4063
rect 6920 4020 6972 4029
rect 7748 4088 7800 4140
rect 10876 4156 10928 4208
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 6552 3884 6604 3936
rect 7104 3884 7156 3936
rect 9036 3952 9088 4004
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9864 4020 9916 4072
rect 10784 4088 10836 4140
rect 10232 3952 10284 4004
rect 7748 3884 7800 3936
rect 8576 3884 8628 3936
rect 9588 3884 9640 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 2412 3680 2464 3732
rect 1676 3587 1728 3596
rect 1676 3553 1685 3587
rect 1685 3553 1719 3587
rect 1719 3553 1728 3587
rect 1676 3544 1728 3553
rect 2412 3544 2464 3596
rect 7288 3587 7340 3596
rect 7288 3553 7297 3587
rect 7297 3553 7331 3587
rect 7331 3553 7340 3587
rect 7288 3544 7340 3553
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 9312 3587 9364 3596
rect 9312 3553 9321 3587
rect 9321 3553 9355 3587
rect 9355 3553 9364 3587
rect 9312 3544 9364 3553
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 10232 3544 10284 3596
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 7840 3519 7892 3528
rect 7840 3485 7849 3519
rect 7849 3485 7883 3519
rect 7883 3485 7892 3519
rect 7840 3476 7892 3485
rect 3976 3408 4028 3460
rect 5540 3451 5592 3460
rect 5540 3417 5549 3451
rect 5549 3417 5583 3451
rect 5583 3417 5592 3451
rect 5540 3408 5592 3417
rect 7196 3408 7248 3460
rect 10600 3408 10652 3460
rect 7380 3383 7432 3392
rect 7380 3349 7389 3383
rect 7389 3349 7423 3383
rect 7423 3349 7432 3383
rect 7380 3340 7432 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5540 3136 5592 3188
rect 7196 3179 7248 3188
rect 2596 3068 2648 3120
rect 3976 3068 4028 3120
rect 7196 3145 7205 3179
rect 7205 3145 7239 3179
rect 7239 3145 7248 3179
rect 7196 3136 7248 3145
rect 7380 3068 7432 3120
rect 8576 3111 8628 3120
rect 8576 3077 8585 3111
rect 8585 3077 8619 3111
rect 8619 3077 8628 3111
rect 8576 3068 8628 3077
rect 9956 3136 10008 3188
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 13268 3068 13320 3120
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 6368 2932 6420 2984
rect 6920 3000 6972 3052
rect 7288 3000 7340 3052
rect 10324 3000 10376 3052
rect 8208 2932 8260 2984
rect 9312 2932 9364 2984
rect 10140 2932 10192 2984
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 7196 2456 7248 2508
rect 7748 2388 7800 2440
rect 7840 2388 7892 2440
rect 7104 2252 7156 2304
rect 7748 2252 7800 2304
rect 8392 2252 8444 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 5814 16333 5870 17133
rect 6458 16333 6514 17133
rect 7102 16333 7158 17133
rect 8390 16333 8446 17133
rect 9678 16333 9734 17133
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 5828 14482 5856 16333
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 6368 14408 6420 14414
rect 6472 14396 6500 16333
rect 7116 14414 7144 16333
rect 8404 14414 8432 16333
rect 9692 14618 9720 16333
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 6420 14368 6500 14396
rect 7104 14408 7156 14414
rect 6368 14350 6420 14356
rect 7104 14350 7156 14356
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 5816 14272 5868 14278
rect 5816 14214 5868 14220
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 5460 13530 5488 13806
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 13161 888 13262
rect 1584 13184 1636 13190
rect 846 13152 902 13161
rect 1584 13126 1636 13132
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 846 13087 902 13096
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1412 11898 1440 12242
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 940 11688 992 11694
rect 938 11656 940 11665
rect 992 11656 994 11665
rect 938 11591 994 11600
rect 1412 10130 1440 11834
rect 1596 11830 1624 13126
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2700 12306 2728 12922
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 2884 12306 2912 12718
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2872 12300 2924 12306
rect 2872 12242 2924 12248
rect 1768 12232 1820 12238
rect 1768 12174 1820 12180
rect 1780 11898 1808 12174
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2608 11898 2636 12038
rect 1768 11892 1820 11898
rect 1768 11834 1820 11840
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2700 11830 2728 12242
rect 2964 12164 3016 12170
rect 2964 12106 3016 12112
rect 1584 11824 1636 11830
rect 1584 11766 1636 11772
rect 2688 11824 2740 11830
rect 2688 11766 2740 11772
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 1952 11552 2004 11558
rect 1952 11494 2004 11500
rect 1964 11150 1992 11494
rect 2516 11150 2544 11698
rect 2976 11694 3004 12106
rect 2964 11688 3016 11694
rect 2700 11648 2964 11676
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 2504 11144 2556 11150
rect 2504 11086 2556 11092
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 846 9072 902 9081
rect 846 9007 902 9016
rect 860 8974 888 9007
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 1688 8634 1716 9454
rect 1872 9178 1900 9930
rect 2228 9512 2280 9518
rect 2228 9454 2280 9460
rect 2240 9382 2268 9454
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1780 8498 1808 8910
rect 2136 8832 2188 8838
rect 2136 8774 2188 8780
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1412 8265 1440 8434
rect 1398 8256 1454 8265
rect 1398 8191 1454 8200
rect 2148 7886 2176 8774
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 938 7576 994 7585
rect 938 7511 994 7520
rect 848 6792 900 6798
rect 846 6760 848 6769
rect 900 6760 902 6769
rect 846 6695 902 6704
rect 952 6322 980 7511
rect 1872 7410 1900 7686
rect 2056 7478 2084 7822
rect 2044 7472 2096 7478
rect 2044 7414 2096 7420
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1688 6390 1716 7346
rect 2056 6866 2084 7414
rect 2240 6914 2268 9318
rect 2320 9104 2372 9110
rect 2320 9046 2372 9052
rect 2332 7392 2360 9046
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2424 8566 2452 8774
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2516 7546 2544 11086
rect 2700 9042 2728 11648
rect 2964 11630 3016 11636
rect 3252 11354 3280 12718
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3528 11286 3556 12174
rect 3712 12170 3740 12378
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 9586 3280 11154
rect 3712 10062 3740 12106
rect 3804 10146 3832 12854
rect 3896 12424 3924 13126
rect 4632 12646 4660 13330
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3896 12396 4108 12424
rect 3896 10810 3924 12396
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3988 11286 4016 12242
rect 4080 12238 4108 12396
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4172 11642 4200 12310
rect 4080 11614 4200 11642
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4080 11150 4108 11614
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4632 11082 4660 12582
rect 4724 11694 4752 12718
rect 4816 12306 4844 13398
rect 5460 13326 5488 13466
rect 5552 13326 5580 13738
rect 5632 13456 5684 13462
rect 5632 13398 5684 13404
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4896 12912 4948 12918
rect 4896 12854 4948 12860
rect 4908 12442 4936 12854
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 5000 12374 5028 12786
rect 4988 12368 5040 12374
rect 4988 12310 5040 12316
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4816 11830 4844 12106
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4804 11824 4856 11830
rect 4804 11766 4856 11772
rect 4896 11756 4948 11762
rect 4896 11698 4948 11704
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4724 11354 4752 11494
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4712 11144 4764 11150
rect 4908 11132 4936 11698
rect 4764 11104 4936 11132
rect 4712 11086 4764 11092
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3804 10118 4016 10146
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3528 9178 3556 9454
rect 3516 9172 3568 9178
rect 3516 9114 3568 9120
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2608 8634 2636 8978
rect 2700 8922 2728 8978
rect 2700 8894 2820 8922
rect 3712 8906 3740 9862
rect 3988 9654 4016 10118
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3988 9518 4016 9590
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2792 8362 2820 8894
rect 3700 8900 3752 8906
rect 3700 8842 3752 8848
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2780 8356 2832 8362
rect 2780 8298 2832 8304
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2608 7546 2636 7822
rect 2688 7744 2740 7750
rect 2688 7686 2740 7692
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2596 7404 2648 7410
rect 2332 7364 2596 7392
rect 2596 7346 2648 7352
rect 2700 7342 2728 7686
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2240 6886 2452 6914
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1676 6384 1728 6390
rect 1676 6326 1728 6332
rect 940 6316 992 6322
rect 940 6258 992 6264
rect 2424 6254 2452 6886
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2516 6390 2544 6598
rect 2884 6458 2912 8434
rect 2976 7274 3004 8774
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 3068 6866 3096 8774
rect 3712 8498 3740 8842
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3344 7954 3372 8366
rect 3712 8362 3740 8434
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3792 7948 3844 7954
rect 3792 7890 3844 7896
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 3160 6934 3188 7346
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3148 6724 3200 6730
rect 3148 6666 3200 6672
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 2044 6248 2096 6254
rect 2044 6190 2096 6196
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 846 6080 902 6089
rect 846 6015 902 6024
rect 860 5710 888 6015
rect 848 5704 900 5710
rect 848 5646 900 5652
rect 2056 5642 2084 6190
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 2148 5710 2176 6054
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2044 5636 2096 5642
rect 2044 5578 2096 5584
rect 846 5400 902 5409
rect 2056 5370 2084 5578
rect 2148 5370 2176 5646
rect 846 5335 902 5344
rect 2044 5364 2096 5370
rect 860 5234 888 5335
rect 2044 5306 2096 5312
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 2240 5166 2268 5646
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 846 4720 902 4729
rect 846 4655 902 4664
rect 860 4622 888 4655
rect 848 4616 900 4622
rect 848 4558 900 4564
rect 1688 3602 1716 4966
rect 2240 4826 2268 5102
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2320 4072 2372 4078
rect 2424 4060 2452 6190
rect 2504 6112 2556 6118
rect 2504 6054 2556 6060
rect 2516 4622 2544 6054
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2516 4214 2544 4422
rect 2504 4208 2556 4214
rect 2504 4150 2556 4156
rect 2372 4032 2452 4060
rect 2320 4014 2372 4020
rect 2424 3738 2452 4032
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2424 3602 2452 3674
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2424 3058 2452 3538
rect 2608 3126 2636 4966
rect 2976 4690 3004 5578
rect 3068 5370 3096 5714
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3160 5166 3188 6666
rect 3252 5914 3280 7142
rect 3344 6798 3372 7686
rect 3804 7410 3832 7890
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3608 7404 3660 7410
rect 3608 7346 3660 7352
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3620 7002 3648 7346
rect 3608 6996 3660 7002
rect 3608 6938 3660 6944
rect 3896 6798 3924 7414
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 5914 3648 6598
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3608 5908 3660 5914
rect 3608 5850 3660 5856
rect 3804 5846 3832 6734
rect 3988 6254 4016 9454
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9058 4660 10746
rect 4724 9110 4752 11086
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4540 9030 4660 9058
rect 4712 9104 4764 9110
rect 4712 9046 4764 9052
rect 4356 8906 4384 8978
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4540 8362 4568 9030
rect 4816 8974 4844 9318
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4080 7818 4108 8230
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7954 4660 8910
rect 4436 7948 4488 7954
rect 4436 7890 4488 7896
rect 4620 7948 4672 7954
rect 4620 7890 4672 7896
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 4448 7410 4476 7890
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4436 7404 4488 7410
rect 4436 7346 4488 7352
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4172 6390 4200 6666
rect 4356 6458 4384 6802
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 4724 6322 4752 7754
rect 4816 7732 4844 8910
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5080 8288 5132 8294
rect 5080 8230 5132 8236
rect 5092 8090 5120 8230
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 4896 7744 4948 7750
rect 4816 7704 4896 7732
rect 4896 7686 4948 7692
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7478 5304 13194
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12850 5488 13126
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5368 12730 5396 12786
rect 5552 12730 5580 13262
rect 5644 12986 5672 13398
rect 5828 13394 5856 14214
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5920 13530 5948 13670
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5816 13388 5868 13394
rect 5816 13330 5868 13336
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5632 12980 5684 12986
rect 5632 12922 5684 12928
rect 5736 12918 5764 13262
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5828 12782 5856 13330
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5724 12776 5776 12782
rect 5368 12702 5488 12730
rect 5552 12724 5724 12730
rect 5552 12718 5776 12724
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 5552 12702 5764 12718
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5368 11694 5396 12378
rect 5460 11762 5488 12702
rect 5920 12306 5948 13126
rect 6104 12986 6132 14282
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 6840 13870 6868 14214
rect 7852 14006 7880 14214
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6380 12850 6408 13194
rect 6644 12912 6696 12918
rect 6644 12854 6696 12860
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 6000 12164 6052 12170
rect 6000 12106 6052 12112
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 11218 5580 11494
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 9518 5580 11018
rect 5736 10810 5764 11698
rect 6012 11082 6040 12106
rect 6472 11626 6500 12650
rect 6552 12096 6604 12102
rect 6656 12084 6684 12854
rect 6932 12714 6960 13670
rect 7024 13530 7052 13874
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6932 12306 6960 12650
rect 7024 12442 7052 12786
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 7116 12186 7144 12582
rect 6604 12056 6684 12084
rect 7024 12158 7144 12186
rect 6552 12038 6604 12044
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6932 11762 6960 11834
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7024 11694 7052 12158
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7116 11694 7144 12038
rect 7208 11898 7236 13670
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7300 12374 7328 13466
rect 7852 13326 7880 13942
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7576 12434 7604 13194
rect 8036 12918 8064 14010
rect 8484 13796 8536 13802
rect 8484 13738 8536 13744
rect 8496 12986 8524 13738
rect 8680 13326 8708 14214
rect 10336 14074 10364 14350
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 9404 13932 9456 13938
rect 9404 13874 9456 13880
rect 9772 13932 9824 13938
rect 9772 13874 9824 13880
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8680 12918 8708 13262
rect 8024 12912 8076 12918
rect 8024 12854 8076 12860
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7484 12406 7604 12434
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 7116 10810 7144 11630
rect 7208 11150 7236 11834
rect 7484 11830 7512 12406
rect 7944 12170 7972 12786
rect 8036 12238 8064 12854
rect 8668 12776 8720 12782
rect 8772 12730 8800 13670
rect 9416 13462 9444 13874
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 8852 13184 8904 13190
rect 8852 13126 8904 13132
rect 8864 12850 8892 13126
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8720 12724 8800 12730
rect 8668 12718 8800 12724
rect 8680 12702 8800 12718
rect 9416 12646 9444 13398
rect 9784 12986 9812 13874
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9968 12714 9996 13806
rect 10704 13394 10732 13874
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10508 13252 10560 13258
rect 10508 13194 10560 13200
rect 10520 12918 10548 13194
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10048 12776 10100 12782
rect 10048 12718 10100 12724
rect 9956 12708 10008 12714
rect 9956 12650 10008 12656
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7564 12164 7616 12170
rect 7564 12106 7616 12112
rect 7932 12164 7984 12170
rect 7932 12106 7984 12112
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7576 11762 7604 12106
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7840 11756 7892 11762
rect 7840 11698 7892 11704
rect 7564 11552 7616 11558
rect 7564 11494 7616 11500
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 6368 10736 6420 10742
rect 6368 10678 6420 10684
rect 6380 9722 6408 10678
rect 7576 10674 7604 11494
rect 7852 11082 7880 11698
rect 8036 11150 8064 12174
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 8576 10600 8628 10606
rect 8576 10542 8628 10548
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8838 5396 8910
rect 5552 8838 5580 9318
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5368 8430 5396 8774
rect 5356 8424 5408 8430
rect 5408 8384 5488 8412
rect 5356 8366 5408 8372
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5368 7818 5396 8026
rect 5460 7886 5488 8384
rect 5552 7886 5580 8774
rect 5644 8634 5672 9114
rect 5828 9110 5856 9454
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5644 8294 5672 8570
rect 5736 8498 5764 8978
rect 5920 8974 5948 9318
rect 6104 9178 6132 9522
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5908 8968 5960 8974
rect 5960 8928 6040 8956
rect 5908 8910 5960 8916
rect 6012 8514 6040 8928
rect 6104 8634 6132 9114
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 5724 8492 5776 8498
rect 6012 8486 6132 8514
rect 5724 8434 5776 8440
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5736 8090 5764 8434
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5356 7812 5408 7818
rect 5356 7754 5408 7760
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 5368 7342 5396 7754
rect 5460 7410 5488 7822
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5356 7336 5408 7342
rect 5356 7278 5408 7284
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5368 6458 5396 7278
rect 5644 6914 5672 7890
rect 5460 6886 5672 6914
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5460 6390 5488 6886
rect 5828 6390 5856 8298
rect 6104 7954 6132 8486
rect 6196 8362 6224 9046
rect 6288 9042 6316 9522
rect 6472 9178 6500 9522
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 8838 6316 8978
rect 6368 8900 6420 8906
rect 6368 8842 6420 8848
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6380 8566 6408 8842
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6472 8498 6500 8774
rect 6564 8634 6592 9590
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6840 9178 6868 9522
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6736 9036 6788 9042
rect 6788 8996 6868 9024
rect 6736 8978 6788 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6460 8492 6512 8498
rect 6460 8434 6512 8440
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6472 8022 6500 8434
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6380 7478 6408 7686
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3160 4690 3188 5102
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3436 3534 3464 4762
rect 3988 4214 4016 6190
rect 4816 6186 4844 6258
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4816 5710 4844 6122
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 5368 5574 5396 6258
rect 5448 6248 5500 6254
rect 5540 6248 5592 6254
rect 5500 6208 5540 6236
rect 5448 6190 5500 6196
rect 5540 6190 5592 6196
rect 5460 5642 5488 6190
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5448 5636 5500 5642
rect 5448 5578 5500 5584
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 4816 5234 4844 5510
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 5368 5166 5396 5510
rect 5460 5234 5488 5578
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 5000 4622 5028 4966
rect 4988 4616 5040 4622
rect 4988 4558 5040 4564
rect 5368 4554 5396 5102
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 5460 4214 5488 5170
rect 5552 5098 5580 6054
rect 5736 5846 5764 6258
rect 6196 5846 6224 7346
rect 6472 6322 6500 7958
rect 6564 7886 6592 8570
rect 6656 8498 6684 8910
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6748 8294 6776 8842
rect 6840 8838 6868 8996
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6564 6254 6592 7822
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 7478 6868 7754
rect 6932 7546 6960 10542
rect 8588 10062 8616 10542
rect 9048 10266 9076 11154
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9036 10260 9088 10266
rect 9036 10202 9088 10208
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7932 9580 7984 9586
rect 7932 9522 7984 9528
rect 7024 8634 7052 9522
rect 7944 8974 7972 9522
rect 8312 9518 8340 9998
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 8128 8838 8156 9318
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 8128 8498 8156 8774
rect 8220 8566 8248 8842
rect 8312 8634 8340 9454
rect 8404 9042 8432 9862
rect 8588 9654 8616 9998
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8772 9722 8800 9862
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 8560 8260 8566
rect 8208 8502 8260 8508
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8220 8430 8248 8502
rect 8208 8424 8260 8430
rect 8312 8401 8340 8570
rect 8588 8430 8616 9590
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8772 9178 8800 9454
rect 8760 9172 8812 9178
rect 8760 9114 8812 9120
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8576 8424 8628 8430
rect 8208 8366 8260 8372
rect 8298 8392 8354 8401
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6748 5914 6776 6258
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 5736 5234 5764 5782
rect 5908 5772 5960 5778
rect 5908 5714 5960 5720
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5552 4758 5580 5034
rect 5736 4826 5764 5170
rect 5920 4826 5948 5714
rect 6840 5710 6868 6394
rect 7116 6322 7144 7346
rect 8220 6798 8248 8366
rect 8576 8366 8628 8372
rect 8298 8327 8354 8336
rect 8588 7886 8616 8366
rect 8680 8294 8708 8978
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8772 8498 8800 8910
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8758 8392 8814 8401
rect 8758 8327 8814 8336
rect 8772 8294 8800 8327
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8864 8022 8892 8910
rect 8956 8906 8984 9046
rect 8944 8900 8996 8906
rect 8944 8842 8996 8848
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8852 8016 8904 8022
rect 8852 7958 8904 7964
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 8116 6316 8168 6322
rect 8116 6258 8168 6264
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6644 5704 6696 5710
rect 6644 5646 6696 5652
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 5724 4820 5776 4826
rect 5724 4762 5776 4768
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5540 4752 5592 4758
rect 5540 4694 5592 4700
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 5448 4208 5500 4214
rect 5448 4150 5500 4156
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3988 3466 4016 4150
rect 5552 4078 5580 4694
rect 6012 4622 6040 5238
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6104 4826 6132 5170
rect 6288 5166 6316 5646
rect 6472 5302 6500 5646
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 6564 5234 6592 5510
rect 6552 5228 6604 5234
rect 6552 5170 6604 5176
rect 6276 5160 6328 5166
rect 6276 5102 6328 5108
rect 6092 4820 6144 4826
rect 6092 4762 6144 4768
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5828 4146 5856 4490
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 5540 3460 5592 3466
rect 5540 3402 5592 3408
rect 3988 3126 4016 3402
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5552 3194 5580 3402
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 6380 2990 6408 4558
rect 6656 4554 6684 5646
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6932 4078 6960 6258
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 7024 5370 7052 6190
rect 8024 6180 8076 6186
rect 8024 6122 8076 6128
rect 8036 5710 8064 6122
rect 8128 5710 8156 6258
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 5574 8156 5646
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 8220 5166 8248 5782
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 7012 4548 7064 4554
rect 7012 4490 7064 4496
rect 7024 4146 7052 4490
rect 7300 4146 7328 5102
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 7852 4214 7880 4626
rect 8312 4554 8340 6258
rect 8404 5710 8432 6258
rect 8496 5778 8524 6802
rect 8772 6390 8800 7482
rect 8864 7342 8892 7958
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8852 6928 8904 6934
rect 8852 6870 8904 6876
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8864 5846 8892 6870
rect 8956 6458 8984 8570
rect 9048 6866 9076 9862
rect 9140 8974 9168 10610
rect 9232 10062 9260 11834
rect 9416 11830 9444 12582
rect 10060 12442 10088 12718
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9508 11898 9536 12174
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9404 11824 9456 11830
rect 9404 11766 9456 11772
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9324 11354 9352 11630
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9416 11121 9444 11766
rect 9508 11150 9536 11834
rect 9496 11144 9548 11150
rect 9402 11112 9458 11121
rect 9496 11086 9548 11092
rect 9402 11047 9458 11056
rect 9600 10826 9628 12242
rect 10244 12238 10272 12786
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10416 11756 10468 11762
rect 10520 11744 10548 12854
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11808 12374 11836 12718
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10468 11716 10548 11744
rect 10416 11698 10468 11704
rect 9416 10798 9628 10826
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 9324 9722 9352 9862
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9128 8968 9180 8974
rect 9416 8922 9444 10798
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9722 9536 9930
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9600 9654 9628 10610
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 9654 9996 10406
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9600 9042 9628 9590
rect 10336 9586 10364 9862
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9128 8910 9180 8916
rect 9140 8634 9168 8910
rect 9324 8894 9444 8922
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9220 8424 9272 8430
rect 9218 8392 9220 8401
rect 9272 8392 9274 8401
rect 9218 8327 9274 8336
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 7546 9260 7822
rect 9324 7546 9352 8894
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 8498 9444 8774
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9220 7540 9272 7546
rect 9220 7482 9272 7488
rect 9312 7540 9364 7546
rect 9312 7482 9364 7488
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 5914 8984 6190
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8496 5098 8524 5714
rect 8852 5704 8904 5710
rect 8852 5646 8904 5652
rect 8484 5092 8536 5098
rect 8484 5034 8536 5040
rect 8864 4622 8892 5646
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8220 4282 8340 4298
rect 8220 4276 8352 4282
rect 8220 4270 8300 4276
rect 7840 4208 7892 4214
rect 7840 4150 7892 4156
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6552 3936 6604 3942
rect 7104 3936 7156 3942
rect 6552 3878 6604 3884
rect 6932 3884 7104 3890
rect 6932 3878 7156 3884
rect 6564 3058 6592 3878
rect 6932 3862 7144 3878
rect 6932 3058 6960 3862
rect 7300 3602 7328 4082
rect 7760 3942 7788 4082
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7196 3460 7248 3466
rect 7196 3402 7248 3408
rect 7208 3194 7236 3402
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7300 3058 7328 3538
rect 7760 3534 7788 3878
rect 7852 3534 7880 4150
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 3126 7420 3334
rect 7380 3120 7432 3126
rect 7380 3062 7432 3068
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 7300 2774 7328 2994
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7208 2746 7328 2774
rect 7208 2514 7236 2746
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 7760 2446 7788 3470
rect 7852 2446 7880 3470
rect 8220 2990 8248 4270
rect 8300 4218 8352 4224
rect 9048 4010 9076 6258
rect 9140 5846 9168 7346
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6254 9260 6734
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9324 5914 9352 7346
rect 9416 7324 9444 8434
rect 9600 7886 9628 8978
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7478 9536 7686
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9876 7410 9904 9454
rect 10060 9178 10088 9454
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 9416 7296 9628 7324
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 6458 9444 6598
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9508 6254 9536 7142
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 9220 5636 9272 5642
rect 9220 5578 9272 5584
rect 9232 5522 9260 5578
rect 9404 5568 9456 5574
rect 9232 5516 9404 5522
rect 9232 5510 9456 5516
rect 9232 5494 9444 5510
rect 9232 4554 9260 5494
rect 9508 4826 9536 6190
rect 9600 6186 9628 7296
rect 9784 6866 9812 7346
rect 10244 6934 10272 7346
rect 10232 6928 10284 6934
rect 10232 6870 10284 6876
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9692 6118 9720 6734
rect 10152 6186 10180 6734
rect 10416 6656 10468 6662
rect 10416 6598 10468 6604
rect 10428 6390 10456 6598
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 10336 5710 10364 6258
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9496 4820 9548 4826
rect 9496 4762 9548 4768
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9232 4078 9260 4490
rect 9876 4282 9904 5510
rect 10060 5234 10088 5578
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10060 4282 10088 5170
rect 10244 5098 10272 5510
rect 10336 5166 10364 5646
rect 10324 5160 10376 5166
rect 10324 5102 10376 5108
rect 10232 5092 10284 5098
rect 10232 5034 10284 5040
rect 10244 4622 10272 5034
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9876 4078 9904 4218
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9036 4004 9088 4010
rect 9036 3946 9088 3952
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 8588 3126 8616 3878
rect 9310 3632 9366 3641
rect 9600 3602 9628 3878
rect 9310 3567 9312 3576
rect 9364 3567 9366 3576
rect 9588 3596 9640 3602
rect 9312 3538 9364 3544
rect 9588 3538 9640 3544
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 9324 2990 9352 3538
rect 9968 3194 9996 4082
rect 10060 3584 10088 4218
rect 10244 4010 10272 4558
rect 10232 4004 10284 4010
rect 10232 3946 10284 3952
rect 10244 3602 10272 3946
rect 10232 3596 10284 3602
rect 10060 3556 10180 3584
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10152 2990 10180 3556
rect 10232 3538 10284 3544
rect 10244 3040 10272 3538
rect 10520 3482 10548 11716
rect 10888 9654 10916 12242
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11164 10674 11192 11222
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11440 10470 11468 11086
rect 11704 11076 11756 11082
rect 11704 11018 11756 11024
rect 12716 11076 12768 11082
rect 12716 11018 12768 11024
rect 13176 11076 13228 11082
rect 13176 11018 13228 11024
rect 11716 10810 11744 11018
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11900 10674 11928 10950
rect 11888 10668 11940 10674
rect 11888 10610 11940 10616
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11428 10464 11480 10470
rect 11428 10406 11480 10412
rect 11440 10062 11468 10406
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 10876 9648 10928 9654
rect 10876 9590 10928 9596
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10692 9580 10744 9586
rect 10692 9522 10744 9528
rect 10612 7546 10640 9522
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10704 6458 10732 9522
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11072 7954 11100 8502
rect 11164 8294 11192 8910
rect 11256 8430 11284 9114
rect 11440 8430 11468 9998
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11716 9722 11744 9930
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11808 9586 11836 10542
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 9586 11928 10474
rect 12268 9738 12296 10610
rect 12440 10600 12492 10606
rect 12360 10548 12440 10554
rect 12360 10542 12492 10548
rect 12360 10526 12480 10542
rect 12360 10470 12388 10526
rect 12348 10464 12400 10470
rect 12348 10406 12400 10412
rect 12728 9994 12756 11018
rect 13188 10742 13216 11018
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 12176 9722 12296 9738
rect 12164 9716 12296 9722
rect 12216 9710 12296 9716
rect 12164 9658 12216 9664
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 8650 11928 9522
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12176 9178 12204 9454
rect 12164 9172 12216 9178
rect 12164 9114 12216 9120
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11716 8622 11928 8650
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11164 8090 11192 8230
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11164 7818 11192 8026
rect 11256 7886 11284 8366
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11152 7812 11204 7818
rect 11152 7754 11204 7760
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10692 6112 10744 6118
rect 10692 6054 10744 6060
rect 10704 5710 10732 6054
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10704 5302 10732 5646
rect 10796 5642 10824 6394
rect 11072 6390 11100 7686
rect 11440 7342 11468 8366
rect 11716 7868 11744 8622
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11900 8430 11928 8502
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11808 8090 11836 8366
rect 11796 8084 11848 8090
rect 11796 8026 11848 8032
rect 11992 7886 12020 8842
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12084 7886 12112 8774
rect 12268 7886 12296 9710
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12636 8974 12664 9522
rect 12532 8968 12584 8974
rect 12532 8910 12584 8916
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 7886 12480 8774
rect 12544 8430 12572 8910
rect 12636 8634 12664 8910
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12728 8548 12756 9930
rect 13096 9654 13124 9930
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 13096 8974 13124 9590
rect 13188 9586 13216 10678
rect 13358 9616 13414 9625
rect 13176 9580 13228 9586
rect 13358 9551 13414 9560
rect 13176 9522 13228 9528
rect 13372 9450 13400 9551
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13084 8968 13136 8974
rect 13084 8910 13136 8916
rect 13358 8936 13414 8945
rect 13358 8871 13414 8880
rect 13372 8838 13400 8871
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 12808 8560 12860 8566
rect 12728 8520 12808 8548
rect 12860 8520 12940 8548
rect 12808 8502 12860 8508
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12544 8276 12572 8366
rect 12544 8248 12664 8276
rect 11888 7880 11940 7886
rect 11716 7840 11888 7868
rect 11888 7822 11940 7828
rect 11980 7880 12032 7886
rect 11980 7822 12032 7828
rect 12072 7880 12124 7886
rect 12072 7822 12124 7828
rect 12256 7880 12308 7886
rect 12256 7822 12308 7828
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 11900 7732 11928 7822
rect 11900 7704 12112 7732
rect 11428 7336 11480 7342
rect 11428 7278 11480 7284
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10784 5636 10836 5642
rect 10784 5578 10836 5584
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10796 4146 10824 5578
rect 10888 4826 10916 6190
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5710 11100 6054
rect 11440 5778 11468 7278
rect 11900 7002 11928 7278
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 12084 6712 12112 7704
rect 12268 6730 12296 7822
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12360 6866 12388 7686
rect 12452 6866 12480 7822
rect 12636 7818 12664 8248
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12636 6798 12664 7754
rect 12820 7546 12848 7822
rect 12808 7540 12860 7546
rect 12808 7482 12860 7488
rect 12912 7478 12940 8520
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13358 8256 13414 8265
rect 13280 7886 13308 8230
rect 13358 8191 13414 8200
rect 13372 8090 13400 8191
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 7585 13032 7686
rect 12990 7576 13046 7585
rect 12990 7511 13046 7520
rect 12900 7472 12952 7478
rect 12900 7414 12952 7420
rect 12912 6914 12940 7414
rect 12820 6886 12940 6914
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12164 6724 12216 6730
rect 12084 6684 12164 6712
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11152 5704 11204 5710
rect 11152 5646 11204 5652
rect 11164 5370 11192 5646
rect 12084 5574 12112 6684
rect 12164 6666 12216 6672
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12268 6458 12296 6666
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12452 6322 12480 6666
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12452 5914 12480 6258
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12820 5710 12848 6886
rect 12808 5704 12860 5710
rect 12808 5646 12860 5652
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12820 5370 12848 5646
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 13268 5296 13320 5302
rect 13268 5238 13320 5244
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10888 4214 10916 4762
rect 13280 4486 13308 5238
rect 13464 5234 13492 5578
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13372 4865 13400 4966
rect 13358 4856 13414 4865
rect 13358 4791 13414 4800
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10520 3466 10640 3482
rect 10520 3460 10652 3466
rect 10520 3454 10600 3460
rect 10600 3402 10652 3408
rect 10612 3194 10640 3402
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 13280 3126 13308 4422
rect 13464 4185 13492 4558
rect 13450 4176 13506 4185
rect 13450 4111 13506 4120
rect 13268 3120 13320 3126
rect 13268 3062 13320 3068
rect 10324 3052 10376 3058
rect 10244 3012 10324 3040
rect 10324 2994 10376 3000
rect 8208 2984 8260 2990
rect 8208 2926 8260 2932
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 10140 2984 10192 2990
rect 10140 2926 10192 2932
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8392 2304 8444 2310
rect 8392 2246 8444 2252
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 7116 800 7144 2246
rect 7760 800 7788 2246
rect 8404 800 8432 2246
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
<< via2 >>
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 846 13096 902 13152
rect 938 11636 940 11656
rect 940 11636 992 11656
rect 992 11636 994 11656
rect 938 11600 994 11636
rect 846 9016 902 9072
rect 1398 8200 1454 8256
rect 938 7520 994 7576
rect 846 6740 848 6760
rect 848 6740 900 6760
rect 900 6740 902 6760
rect 846 6704 902 6740
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 846 6024 902 6080
rect 846 5344 902 5400
rect 846 4664 902 4720
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 8298 8336 8354 8392
rect 8758 8336 8814 8392
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 9402 11056 9458 11112
rect 9218 8372 9220 8392
rect 9220 8372 9272 8392
rect 9272 8372 9274 8392
rect 9218 8336 9274 8372
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 9310 3596 9366 3632
rect 9310 3576 9312 3596
rect 9312 3576 9364 3596
rect 9364 3576 9366 3596
rect 13358 9560 13414 9616
rect 13358 8880 13414 8936
rect 13358 8200 13414 8256
rect 12990 7520 13046 7576
rect 13358 4800 13414 4856
rect 13450 4120 13506 4176
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 0 12928 800 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 9254 11052 9260 11116
rect 9324 11114 9330 11116
rect 9397 11114 9463 11117
rect 9324 11112 9463 11114
rect 9324 11056 9402 11112
rect 9458 11056 9463 11112
rect 9324 11054 9463 11056
rect 9324 11052 9330 11054
rect 9397 11051 9463 11054
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 13353 9618 13419 9621
rect 14189 9618 14989 9648
rect 13353 9616 14989 9618
rect 13353 9560 13358 9616
rect 13414 9560 14989 9616
rect 13353 9558 14989 9560
rect 13353 9555 13419 9558
rect 14189 9528 14989 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 13353 8938 13419 8941
rect 14189 8938 14989 8968
rect 13353 8936 14989 8938
rect 13353 8880 13358 8936
rect 13414 8880 14989 8936
rect 13353 8878 14989 8880
rect 0 8848 800 8878
rect 13353 8875 13419 8878
rect 14189 8848 14989 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 8293 8394 8359 8397
rect 8753 8394 8819 8397
rect 9213 8394 9279 8397
rect 8293 8392 9279 8394
rect 8293 8336 8298 8392
rect 8354 8336 8758 8392
rect 8814 8336 9218 8392
rect 9274 8336 9279 8392
rect 8293 8334 9279 8336
rect 8293 8331 8359 8334
rect 8753 8331 8819 8334
rect 9213 8331 9279 8334
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 13353 8258 13419 8261
rect 14189 8258 14989 8288
rect 13353 8256 14989 8258
rect 13353 8200 13358 8256
rect 13414 8200 14989 8256
rect 13353 8198 14989 8200
rect 13353 8195 13419 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 14189 8168 14989 8198
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 933 7578 999 7581
rect 0 7576 999 7578
rect 0 7520 938 7576
rect 994 7520 999 7576
rect 0 7518 999 7520
rect 0 7488 800 7518
rect 933 7515 999 7518
rect 12985 7578 13051 7581
rect 14189 7578 14989 7608
rect 12985 7576 14989 7578
rect 12985 7520 12990 7576
rect 13046 7520 14989 7576
rect 12985 7518 14989 7520
rect 12985 7515 13051 7518
rect 14189 7488 14989 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 0 6808 858 6898
rect 798 6765 858 6808
rect 798 6760 907 6765
rect 798 6704 846 6760
rect 902 6704 907 6760
rect 798 6702 907 6704
rect 841 6699 907 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6218 800 6248
rect 0 6128 858 6218
rect 798 6085 858 6128
rect 798 6080 907 6085
rect 798 6024 846 6080
rect 902 6024 907 6080
rect 798 6022 907 6024
rect 841 6019 907 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 0 5538 800 5568
rect 0 5448 858 5538
rect 798 5405 858 5448
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 798 5400 907 5405
rect 798 5344 846 5400
rect 902 5344 907 5400
rect 798 5342 907 5344
rect 841 5339 907 5342
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 13353 4858 13419 4861
rect 14189 4858 14989 4888
rect 0 4768 858 4858
rect 13353 4856 14989 4858
rect 13353 4800 13358 4856
rect 13414 4800 14989 4856
rect 13353 4798 14989 4800
rect 13353 4795 13419 4798
rect 14189 4768 14989 4798
rect 798 4725 858 4768
rect 798 4720 907 4725
rect 798 4664 846 4720
rect 902 4664 907 4720
rect 798 4662 907 4664
rect 841 4659 907 4662
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 13445 4178 13511 4181
rect 14189 4178 14989 4208
rect 13445 4176 14989 4178
rect 13445 4120 13450 4176
rect 13506 4120 14989 4176
rect 13445 4118 14989 4120
rect 13445 4115 13511 4118
rect 14189 4088 14989 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 9305 3636 9371 3637
rect 9254 3572 9260 3636
rect 9324 3634 9371 3636
rect 9324 3632 9416 3634
rect 9366 3576 9416 3632
rect 9324 3574 9416 3576
rect 9324 3572 9371 3574
rect 9305 3571 9371 3572
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 9260 11052 9324 11116
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 9260 3632 9324 3636
rect 9260 3576 9310 3632
rect 9310 3576 9324 3632
rect 9260 3572 9324 3576
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 14720 4528 14736
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 14176 5188 14736
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 9259 11116 9325 11117
rect 9259 11052 9260 11116
rect 9324 11052 9325 11116
rect 9259 11051 9325 11052
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 9262 3637 9322 11051
rect 9259 3636 9325 3637
rect 9259 3572 9260 3636
rect 9324 3572 9325 3636
rect 9259 3571 9325 3572
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _140_
timestamp -25199
transform 1 0 7912 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp -25199
transform -1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp -25199
transform 1 0 8740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _143_
timestamp -25199
transform 1 0 8096 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _144_
timestamp -25199
transform -1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _145_
timestamp -25199
transform 1 0 7544 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _146_
timestamp -25199
transform 1 0 8004 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _147_
timestamp -25199
transform -1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _148_
timestamp -25199
transform -1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _149_
timestamp -25199
transform 1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _150_
timestamp -25199
transform -1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _151_
timestamp -25199
transform 1 0 9476 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _152_
timestamp -25199
transform 1 0 8188 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _153_
timestamp -25199
transform -1 0 8832 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _154_
timestamp -25199
transform 1 0 8004 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _155_
timestamp -25199
transform -1 0 9476 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _156_
timestamp -25199
transform 1 0 8188 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _157_
timestamp -25199
transform 1 0 8924 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _158_
timestamp -25199
transform -1 0 10028 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _159_
timestamp -25199
transform 1 0 8740 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _160_
timestamp -25199
transform 1 0 8188 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _161_
timestamp -25199
transform -1 0 7636 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _162_
timestamp -25199
transform -1 0 8096 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _163_
timestamp -25199
transform -1 0 6992 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp -25199
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _165_
timestamp -25199
transform 1 0 6716 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _166_
timestamp -25199
transform 1 0 7636 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _167_
timestamp -25199
transform 1 0 6716 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _168_
timestamp -25199
transform 1 0 9752 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _169_
timestamp -25199
transform 1 0 5612 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _170_
timestamp -25199
transform 1 0 7452 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _171_
timestamp -25199
transform -1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _172_
timestamp -25199
transform 1 0 8740 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _173_
timestamp -25199
transform -1 0 10396 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _174_
timestamp -25199
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _175_
timestamp -25199
transform -1 0 9568 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _176_
timestamp -25199
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _177_
timestamp -25199
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _178_
timestamp -25199
transform -1 0 2484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_4  _179_
timestamp -25199
transform -1 0 2944 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_2  _180_
timestamp -25199
transform 1 0 2208 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _181_
timestamp -25199
transform 1 0 1656 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _182_
timestamp -25199
transform -1 0 5060 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _183_
timestamp -25199
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _184_
timestamp -25199
transform 1 0 2944 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _185_
timestamp -25199
transform -1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _186_
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _187_
timestamp -25199
transform 1 0 2668 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _188_
timestamp -25199
transform -1 0 4416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _189_
timestamp -25199
transform -1 0 3956 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _190_
timestamp -25199
transform -1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _191_
timestamp -25199
transform -1 0 4876 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _192_
timestamp -25199
transform -1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _193_
timestamp -25199
transform 1 0 2116 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _194_
timestamp -25199
transform 1 0 3588 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _195_
timestamp -25199
transform 1 0 3772 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_2  _196_
timestamp -25199
transform -1 0 4784 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _197_
timestamp -25199
transform -1 0 6072 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _198_
timestamp -25199
transform -1 0 8648 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _199_
timestamp -25199
transform 1 0 9292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _200_
timestamp -25199
transform -1 0 10396 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp -25199
transform 1 0 9108 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _202_
timestamp -25199
transform -1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _203_
timestamp -25199
transform 1 0 7820 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _204_
timestamp -25199
transform -1 0 5336 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _205_
timestamp -25199
transform 1 0 5428 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _206_
timestamp -25199
transform 1 0 9936 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _207_
timestamp -25199
transform 1 0 8372 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _208_
timestamp -25199
transform 1 0 5336 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _209_
timestamp -25199
transform -1 0 5704 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _210_
timestamp -25199
transform 1 0 5796 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _211_
timestamp -25199
transform -1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _212_
timestamp -25199
transform 1 0 5888 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _213_
timestamp -25199
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _214_
timestamp -25199
transform 1 0 4968 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _215_
timestamp -25199
transform -1 0 6348 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _216_
timestamp -25199
transform -1 0 6992 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _217_
timestamp -25199
transform 1 0 5152 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _218_
timestamp -25199
transform 1 0 5612 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _219_
timestamp -25199
transform 1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _220_
timestamp -25199
transform -1 0 6532 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _221_
timestamp -25199
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _222_
timestamp -25199
transform 1 0 6256 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _223_
timestamp -25199
transform 1 0 4784 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _224_
timestamp -25199
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _225_
timestamp -25199
transform 1 0 6348 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _226_
timestamp -25199
transform 1 0 4968 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _227_
timestamp -25199
transform 1 0 5612 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _228_
timestamp -25199
transform 1 0 5612 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _229_
timestamp -25199
transform -1 0 7176 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o31ai_1  _230_
timestamp -25199
transform 1 0 5336 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _231_
timestamp -25199
transform -1 0 7084 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp -25199
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _233_
timestamp -25199
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _234_
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _235_
timestamp -25199
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _236_
timestamp -25199
transform 1 0 5704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp -25199
transform -1 0 10304 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _238_
timestamp -25199
transform -1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _239_
timestamp -25199
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a221oi_1  _240_
timestamp -25199
transform -1 0 9476 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _241_
timestamp -25199
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _242_
timestamp -25199
transform 1 0 9476 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _243_
timestamp -25199
transform 1 0 10212 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _244_
timestamp -25199
transform -1 0 11316 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _245_
timestamp -25199
transform -1 0 11132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _246_
timestamp -25199
transform -1 0 10948 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _247_
timestamp -25199
transform 1 0 10028 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _248_
timestamp -25199
transform -1 0 7544 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _249_
timestamp -25199
transform -1 0 7912 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _250_
timestamp -25199
transform -1 0 7820 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp -25199
transform 1 0 8648 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _252_
timestamp -25199
transform -1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _253_
timestamp -25199
transform 1 0 9752 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _254_
timestamp -25199
transform 1 0 7360 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _255_
timestamp -25199
transform -1 0 7360 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _256_
timestamp -25199
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _257_
timestamp -25199
transform 1 0 10028 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp -25199
transform -1 0 12236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _259_
timestamp -25199
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _260_
timestamp -25199
transform -1 0 11408 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _261_
timestamp -25199
transform 1 0 12512 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _262_
timestamp -25199
transform -1 0 12788 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _263_
timestamp -25199
transform 1 0 11776 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _264_
timestamp -25199
transform 1 0 10948 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp -25199
transform 1 0 12604 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _266_
timestamp -25199
transform 1 0 12052 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _267_
timestamp -25199
transform -1 0 12328 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _268_
timestamp -25199
transform 1 0 12696 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _269_
timestamp -25199
transform -1 0 12696 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _270_
timestamp -25199
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _271_
timestamp -25199
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _272_
timestamp -25199
transform -1 0 12788 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _273_
timestamp -25199
transform -1 0 3588 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _274_
timestamp -25199
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp -25199
transform 1 0 2576 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _276_
timestamp -25199
transform 1 0 2484 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _277_
timestamp -25199
transform 1 0 1748 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp -25199
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _279_
timestamp -25199
transform 1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _280_
timestamp -25199
transform 1 0 2484 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _281_
timestamp -25199
transform 1 0 2024 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _282_
timestamp -25199
transform 1 0 2116 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _283_
timestamp -25199
transform 1 0 4784 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp -25199
transform 1 0 5244 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _285_
timestamp -25199
transform 1 0 5244 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _286_
timestamp -25199
transform -1 0 10764 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _287_
timestamp -25199
transform 1 0 9016 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _288_
timestamp -25199
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _289_
timestamp -25199
transform 1 0 8280 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _290_
timestamp -25199
transform 1 0 9292 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _291_
timestamp -25199
transform 1 0 5244 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _292_
timestamp -25199
transform 1 0 11408 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _293_
timestamp -25199
transform 1 0 11592 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _294_
timestamp -25199
transform 1 0 11500 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _295_
timestamp -25199
transform 1 0 11408 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _296_
timestamp -25199
transform 1 0 11408 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _297_
timestamp -25199
transform 1 0 2852 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _298_
timestamp -25199
transform 1 0 2392 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _299_
timestamp -25199
transform 1 0 2300 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _300_
timestamp -25199
transform 1 0 1380 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _301_
timestamp -25199
transform 1 0 3220 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _302_
timestamp -25199
transform 1 0 1380 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _303_
timestamp -25199
transform 1 0 2484 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _304_
timestamp -25199
transform 1 0 1564 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _305_
timestamp -25199
transform 1 0 1380 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp -25199
transform 1 0 5980 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp -25199
transform 1 0 3036 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxtp_1  _308_
timestamp -25199
transform 1 0 8648 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout24
timestamp -25199
transform 1 0 6992 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout25
timestamp -25199
transform 1 0 4600 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout26
timestamp -25199
transform 1 0 4968 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout27
timestamp -25199
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout28
timestamp -25199
transform -1 0 4140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout29
timestamp -25199
transform -1 0 8648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout30
timestamp -25199
transform -1 0 7636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout31
timestamp -25199
transform -1 0 11040 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout32
timestamp -25199
transform -1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout33
timestamp -25199
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout34
timestamp -25199
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout35
timestamp -25199
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp -25199
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp -25199
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70
timestamp -25199
transform 1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77
timestamp -25199
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636943256
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636943256
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp -25199
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636943256
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_125
timestamp -25199
transform 1 0 12604 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_133
timestamp -25199
transform 1 0 13340 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_3
timestamp -25199
transform 1 0 1380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_11
timestamp -25199
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_34
timestamp 1636943256
transform 1 0 4232 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_46
timestamp -25199
transform 1 0 5336 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp -25199
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_1_71
timestamp -25199
transform 1 0 7636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_77
timestamp -25199
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_98
timestamp -25199
transform 1 0 10120 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp -25199
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636943256
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_125
timestamp -25199
transform 1 0 12604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp -25199
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp -25199
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636943256
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp -25199
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_74
timestamp -25199
transform 1 0 7912 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp -25199
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp -25199
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_112
timestamp 1636943256
transform 1 0 11408 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_124
timestamp -25199
transform 1 0 12512 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_132
timestamp -25199
transform 1 0 13248 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp -25199
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_11
timestamp -25199
transform 1 0 2116 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_36
timestamp 1636943256
transform 1 0 4416 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp -25199
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp -25199
transform 1 0 7360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_76
timestamp -25199
transform 1 0 8096 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_91
timestamp -25199
transform 1 0 9476 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_102
timestamp -25199
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp -25199
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636943256
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_125
timestamp -25199
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp -25199
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp -25199
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp -25199
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636943256
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp -25199
transform 1 0 4876 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_49
timestamp -25199
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_53
timestamp -25199
transform 1 0 5980 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_63
timestamp 1636943256
transform 1 0 6900 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_75
timestamp -25199
transform 1 0 8004 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp -25199
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_92
timestamp -25199
transform 1 0 9568 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_98
timestamp -25199
transform 1 0 10120 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_104
timestamp 1636943256
transform 1 0 10672 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_116
timestamp 1636943256
transform 1 0 11776 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_128
timestamp -25199
transform 1 0 12880 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_6
timestamp -25199
transform 1 0 1656 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_25
timestamp 1636943256
transform 1 0 3404 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_37
timestamp -25199
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_65
timestamp 1636943256
transform 1 0 7084 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_77
timestamp 1636943256
transform 1 0 8188 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_89
timestamp 1636943256
transform 1 0 9292 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_101
timestamp -25199
transform 1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp -25199
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_120
timestamp -25199
transform 1 0 12144 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_130
timestamp -25199
transform 1 0 13064 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp -25199
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp -25199
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636943256
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_41
timestamp -25199
transform 1 0 4876 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_62
timestamp 1636943256
transform 1 0 6808 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_93
timestamp -25199
transform 1 0 9660 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp -25199
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_66
timestamp -25199
transform 1 0 7176 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_82
timestamp -25199
transform 1 0 8648 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_97
timestamp -25199
transform 1 0 10028 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp -25199
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp -25199
transform 1 0 11500 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp -25199
transform 1 0 11868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_121
timestamp 1636943256
transform 1 0 12236 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_133
timestamp -25199
transform 1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp -25199
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_37
timestamp 1636943256
transform 1 0 4508 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_49
timestamp 1636943256
transform 1 0 5612 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_61
timestamp 1636943256
transform 1 0 6716 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_73
timestamp -25199
transform 1 0 7820 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_104
timestamp 1636943256
transform 1 0 10672 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_127
timestamp -25199
transform 1 0 12788 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_9_36
timestamp -25199
transform 1 0 4416 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_64
timestamp 1636943256
transform 1 0 6992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_76
timestamp -25199
transform 1 0 8096 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_100
timestamp 1636943256
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp -25199
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp -25199
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_41
timestamp -25199
transform 1 0 4876 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_64
timestamp 1636943256
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp -25199
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp -25199
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_91
timestamp 1636943256
transform 1 0 9476 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_103
timestamp -25199
transform 1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_34
timestamp 1636943256
transform 1 0 4232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_46
timestamp -25199
transform 1 0 5336 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_50
timestamp -25199
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_61
timestamp 1636943256
transform 1 0 6716 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_73
timestamp -25199
transform 1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_90
timestamp 1636943256
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_102
timestamp -25199
transform 1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_106
timestamp -25199
transform 1 0 10856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_134
timestamp -25199
transform 1 0 13432 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_6
timestamp -25199
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp -25199
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp -25199
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp -25199
transform 1 0 7820 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_101
timestamp 1636943256
transform 1 0 10396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_113
timestamp -25199
transform 1 0 11500 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_128
timestamp -25199
transform 1 0 12880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_43
timestamp -25199
transform 1 0 5060 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_49
timestamp -25199
transform 1 0 5612 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_65
timestamp -25199
transform 1 0 7084 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_73
timestamp -25199
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp -25199
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp -25199
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp -25199
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp -25199
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636943256
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636943256
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1636943256
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1636943256
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_77
timestamp -25199
transform 1 0 8188 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_92
timestamp -25199
transform 1 0 9568 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1636943256
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_109
timestamp -25199
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636943256
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636943256
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636943256
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_39
timestamp -25199
transform 1 0 4692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_47
timestamp -25199
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_57
timestamp -25199
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_73
timestamp 1636943256
transform 1 0 7820 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp -25199
transform 1 0 8924 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_90
timestamp 1636943256
transform 1 0 9384 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_102
timestamp -25199
transform 1 0 10488 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_108
timestamp -25199
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_127
timestamp -25199
transform 1 0 12788 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_3
timestamp -25199
transform 1 0 1380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_11
timestamp -25199
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_17
timestamp -25199
transform 1 0 2668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_25
timestamp -25199
transform 1 0 3404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_35
timestamp -25199
transform 1 0 4324 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_43
timestamp -25199
transform 1 0 5060 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_70
timestamp 1636943256
transform 1 0 7544 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp -25199
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_92
timestamp 1636943256
transform 1 0 9568 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_104
timestamp -25199
transform 1 0 10672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_10
timestamp -25199
transform 1 0 2024 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_20
timestamp -25199
transform 1 0 2944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_41
timestamp -25199
transform 1 0 4876 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_49
timestamp -25199
transform 1 0 5612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_53
timestamp -25199
transform 1 0 5980 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_60
timestamp -25199
transform 1 0 6624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_74
timestamp -25199
transform 1 0 7912 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_82
timestamp -25199
transform 1 0 8648 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_106
timestamp -25199
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636943256
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_125
timestamp -25199
transform 1 0 12604 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp -25199
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp -25199
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_42
timestamp -25199
transform 1 0 4968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp -25199
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_85
timestamp -25199
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_92
timestamp -25199
transform 1 0 9568 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_96
timestamp -25199
transform 1 0 9936 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_104
timestamp 1636943256
transform 1 0 10672 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_116
timestamp 1636943256
transform 1 0 11776 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_128
timestamp -25199
transform 1 0 12880 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp -25199
transform 1 0 13432 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636943256
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_46
timestamp -25199
transform 1 0 5336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp -25199
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_76
timestamp -25199
transform 1 0 8096 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_101
timestamp -25199
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp -25199
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_133
timestamp -25199
transform 1 0 13340 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_6
timestamp 1636943256
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp -25199
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp -25199
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_33
timestamp -25199
transform 1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_78
timestamp -25199
transform 1 0 8280 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_105
timestamp 1636943256
transform 1 0 10764 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_117
timestamp 1636943256
transform 1 0 11868 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_129
timestamp -25199
transform 1 0 12972 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1636943256
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1636943256
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1636943256
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_39
timestamp -25199
transform 1 0 4692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp -25199
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_60
timestamp -25199
transform 1 0 6624 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_67
timestamp 1636943256
transform 1 0 7268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp -25199
transform 1 0 8372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_86
timestamp -25199
transform 1 0 9016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_101
timestamp -25199
transform 1 0 10396 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp -25199
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1636943256
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp -25199
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_133
timestamp -25199
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1636943256
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1636943256
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp -25199
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1636943256
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1636943256
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_69
timestamp -25199
transform 1 0 7452 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_77
timestamp -25199
transform 1 0 8188 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp -25199
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp -25199
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_93
timestamp -25199
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_98
timestamp 1636943256
transform 1 0 10120 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_110
timestamp -25199
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 1636943256
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_125
timestamp -25199
transform 1 0 12604 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp -25199
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp -25199
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -25199
transform -1 0 2024 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp -25199
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  input4
timestamp -25199
transform 1 0 1380 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input5
timestamp -25199
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp -25199
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp -25199
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input8
timestamp -25199
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input9
timestamp -25199
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input10
timestamp -25199
transform -1 0 6256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp -25199
transform -1 0 7452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp -25199
transform 1 0 13248 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp -25199
transform -1 0 8740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output14
timestamp -25199
transform -1 0 10120 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp -25199
transform -1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp -25199
transform -1 0 8188 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp -25199
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp -25199
transform 1 0 13156 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp -25199
transform 1 0 12788 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp -25199
transform 1 0 13156 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp -25199
transform 1 0 13156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp -25199
transform 1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  output23
timestamp -25199
transform 1 0 6348 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_23
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 13800 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_24
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_25
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 13800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_26
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 13800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_27
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 13800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_28
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 13800 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_29
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 13800 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_30
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_31
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 13800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_32
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_33
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 13800 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_34
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 13800 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_35
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 13800 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_36
timestamp -25199
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp -25199
transform -1 0 13800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_37
timestamp -25199
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp -25199
transform -1 0 13800 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_38
timestamp -25199
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp -25199
transform -1 0 13800 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_39
timestamp -25199
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp -25199
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_40
timestamp -25199
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp -25199
transform -1 0 13800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_41
timestamp -25199
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp -25199
transform -1 0 13800 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_42
timestamp -25199
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp -25199
transform -1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_43
timestamp -25199
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp -25199
transform -1 0 13800 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_44
timestamp -25199
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp -25199
transform -1 0 13800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_45
timestamp -25199
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp -25199
transform -1 0 13800 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1
timestamp -25199
transform -1 0 3496 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp -25199
transform -1 0 2116 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer3
timestamp -25199
transform 1 0 2760 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp -25199
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp -25199
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_50
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_51
timestamp -25199
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_52
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_53
timestamp -25199
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_54
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_55
timestamp -25199
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_56
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_57
timestamp -25199
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_58
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_59
timestamp -25199
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_60
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_61
timestamp -25199
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_62
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_63
timestamp -25199
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_64
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_65
timestamp -25199
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_66
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_67
timestamp -25199
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_68
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_69
timestamp -25199
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_70
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_71
timestamp -25199
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_72
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_73
timestamp -25199
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_74
timestamp -25199
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_75
timestamp -25199
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_76
timestamp -25199
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_77
timestamp -25199
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_78
timestamp -25199
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_79
timestamp -25199
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_80
timestamp -25199
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_81
timestamp -25199
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_82
timestamp -25199
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_83
timestamp -25199
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_84
timestamp -25199
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_85
timestamp -25199
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_86
timestamp -25199
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_87
timestamp -25199
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_88
timestamp -25199
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_89
timestamp -25199
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_90
timestamp -25199
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_91
timestamp -25199
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_92
timestamp -25199
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_93
timestamp -25199
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_94
timestamp -25199
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_95
timestamp -25199
transform 1 0 11408 0 1 14144
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 14736 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 14736 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 clk_i
port 2 nsew signal input
flabel metal2 s 9678 16333 9734 17133 0 FreeSans 224 90 0 0 clk_o
port 3 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 cycl_count_o[0]
port 4 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 cycl_count_o[1]
port 5 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 cycl_count_o[2]
port 6 nsew signal output
flabel metal3 s 14189 4768 14989 4888 0 FreeSans 480 0 0 0 cycl_count_o[3]
port 7 nsew signal output
flabel metal3 s 14189 7488 14989 7608 0 FreeSans 480 0 0 0 cycl_count_o[4]
port 8 nsew signal output
flabel metal3 s 14189 8168 14989 8288 0 FreeSans 480 0 0 0 cycl_count_o[5]
port 9 nsew signal output
flabel metal3 s 14189 8848 14989 8968 0 FreeSans 480 0 0 0 cycl_count_o[6]
port 10 nsew signal output
flabel metal3 s 14189 9528 14989 9648 0 FreeSans 480 0 0 0 cycl_count_o[7]
port 11 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 div_i[0]
port 12 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 div_i[1]
port 13 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 div_i[2]
port 14 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 div_i[3]
port 15 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 div_i[4]
port 16 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 div_i[5]
port 17 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 div_i[6]
port 18 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 div_i[7]
port 19 nsew signal input
flabel metal2 s 5814 16333 5870 17133 0 FreeSans 224 90 0 0 div_ready_o
port 20 nsew signal output
flabel metal2 s 6458 16333 6514 17133 0 FreeSans 224 90 0 0 div_valid_i
port 21 nsew signal input
flabel metal2 s 7102 16333 7158 17133 0 FreeSans 224 90 0 0 en_i
port 22 nsew signal input
flabel metal3 s 14189 4088 14989 4208 0 FreeSans 480 0 0 0 rst_ni
port 23 nsew signal input
flabel metal2 s 8390 16333 8446 17133 0 FreeSans 224 90 0 0 test_mode_en_i
port 24 nsew signal input
rlabel metal1 7452 14144 7452 14144 0 VGND
rlabel metal1 7452 14688 7452 14688 0 VPWR
rlabel metal1 8924 12818 8924 12818 0 _000_
rlabel via1 8694 12733 8694 12733 0 _001_
rlabel metal1 10442 13906 10442 13906 0 _002_
rlabel metal1 8970 11662 8970 11662 0 _003_
rlabel metal1 5750 12274 5750 12274 0 _004_
rlabel metal2 5566 11356 5566 11356 0 _005_
rlabel metal1 9430 11322 9430 11322 0 _006_
rlabel metal1 11224 12342 11224 12342 0 _007_
rlabel metal2 8602 3502 8602 3502 0 _008_
rlabel metal2 9614 3740 9614 3740 0 _009_
rlabel metal1 5980 3162 5980 3162 0 _010_
rlabel metal1 11546 5610 11546 5610 0 _011_
rlabel metal1 11868 6970 11868 6970 0 _012_
rlabel metal1 12052 8058 12052 8058 0 _013_
rlabel metal1 11638 9690 11638 9690 0 _014_
rlabel metal1 11960 10778 11960 10778 0 _015_
rlabel metal1 3542 11322 3542 11322 0 _016_
rlabel metal1 2668 3094 2668 3094 0 _017_
rlabel metal1 2576 4182 2576 4182 0 _018_
rlabel metal2 1702 4284 1702 4284 0 _019_
rlabel metal1 3680 9146 3680 9146 0 _020_
rlabel metal1 2116 8602 2116 8602 0 _021_
rlabel metal2 2530 6494 2530 6494 0 _022_
rlabel metal1 1978 9146 1978 9146 0 _023_
rlabel metal1 1978 11866 1978 11866 0 _024_
rlabel metal1 4784 12750 4784 12750 0 _025_
rlabel metal1 9384 6426 9384 6426 0 _026_
rlabel metal1 9568 6698 9568 6698 0 _027_
rlabel metal1 9016 6834 9016 6834 0 _028_
rlabel metal1 9016 10234 9016 10234 0 _029_
rlabel metal1 6118 13770 6118 13770 0 _030_
rlabel metal2 1702 6868 1702 6868 0 _031_
rlabel metal2 2530 9316 2530 9316 0 _032_
rlabel metal1 3726 12206 3726 12206 0 _033_
rlabel metal2 3818 6290 3818 6290 0 _034_
rlabel metal2 4186 6528 4186 6528 0 _035_
rlabel metal1 3542 5882 3542 5882 0 _036_
rlabel via1 3910 6766 3910 6766 0 _037_
rlabel metal1 3772 6698 3772 6698 0 _038_
rlabel metal1 4048 6970 4048 6970 0 _039_
rlabel metal2 3266 6528 3266 6528 0 _040_
rlabel via1 3799 7378 3799 7378 0 _041_
rlabel metal1 2530 7888 2530 7888 0 _042_
rlabel metal2 4094 8024 4094 8024 0 _043_
rlabel metal1 2392 7854 2392 7854 0 _044_
rlabel metal2 2162 8330 2162 8330 0 _045_
rlabel metal2 2714 7514 2714 7514 0 _046_
rlabel metal1 4554 13260 4554 13260 0 _047_
rlabel metal1 4876 13430 4876 13430 0 _048_
rlabel metal1 5566 12818 5566 12818 0 _049_
rlabel metal2 8510 13362 8510 13362 0 _050_
rlabel metal1 9752 12410 9752 12410 0 _051_
rlabel metal2 9798 13430 9798 13430 0 _052_
rlabel metal1 5382 13498 5382 13498 0 _053_
rlabel metal1 5842 9010 5842 9010 0 _054_
rlabel metal1 6210 9146 6210 9146 0 _055_
rlabel metal2 6302 9180 6302 9180 0 _056_
rlabel metal2 6486 9350 6486 9350 0 _057_
rlabel metal1 6762 9520 6762 9520 0 _058_
rlabel metal1 6532 8466 6532 8466 0 _059_
rlabel metal1 6486 7922 6486 7922 0 _060_
rlabel metal2 6394 7582 6394 7582 0 _061_
rlabel metal1 6762 5236 6762 5236 0 _062_
rlabel metal1 6256 5134 6256 5134 0 _063_
rlabel metal2 6578 5372 6578 5372 0 _064_
rlabel metal2 6118 4998 6118 4998 0 _065_
rlabel metal2 7038 5780 7038 5780 0 _066_
rlabel metal1 6578 5882 6578 5882 0 _067_
rlabel metal1 5382 4590 5382 4590 0 _068_
rlabel metal1 5888 4794 5888 4794 0 _069_
rlabel metal2 6946 5168 6946 5168 0 _070_
rlabel metal1 5658 7310 5658 7310 0 _071_
rlabel metal1 6394 7514 6394 7514 0 _072_
rlabel metal2 6210 6596 6210 6596 0 _073_
rlabel metal2 7130 6834 7130 6834 0 _074_
rlabel metal1 6578 8908 6578 8908 0 _075_
rlabel metal1 6946 9146 6946 9146 0 _076_
rlabel metal1 6854 8602 6854 8602 0 _077_
rlabel metal1 6578 10710 6578 10710 0 _078_
rlabel metal2 6946 9044 6946 9044 0 _079_
rlabel metal2 5750 11254 5750 11254 0 _080_
rlabel metal1 9936 7310 9936 7310 0 _081_
rlabel metal1 9338 5814 9338 5814 0 _082_
rlabel metal2 9338 6630 9338 6630 0 _083_
rlabel metal2 9246 7684 9246 7684 0 _084_
rlabel metal2 9522 7582 9522 7582 0 _085_
rlabel metal1 10304 7514 10304 7514 0 _086_
rlabel metal1 10764 4794 10764 4794 0 _087_
rlabel metal2 11086 7038 11086 7038 0 _088_
rlabel metal1 10672 6426 10672 6426 0 _089_
rlabel metal2 10902 10948 10902 10948 0 _090_
rlabel metal1 8418 4046 8418 4046 0 _091_
rlabel metal2 7590 11084 7590 11084 0 _092_
rlabel metal1 12558 10608 12558 10608 0 _093_
rlabel metal1 10120 3162 10120 3162 0 _094_
rlabel metal1 7038 3094 7038 3094 0 _095_
rlabel metal2 6578 3468 6578 3468 0 _096_
rlabel metal2 12466 6086 12466 6086 0 _097_
rlabel metal2 11086 5882 11086 5882 0 _098_
rlabel metal1 11362 5338 11362 5338 0 _099_
rlabel metal1 12098 6664 12098 6664 0 _100_
rlabel metal1 12006 6800 12006 6800 0 _101_
rlabel metal2 12650 8772 12650 8772 0 _102_
rlabel metal2 12006 8364 12006 8364 0 _103_
rlabel metal2 12098 8330 12098 8330 0 _104_
rlabel metal2 11822 10064 11822 10064 0 _105_
rlabel metal1 11730 9452 11730 9452 0 _106_
rlabel metal1 12696 10642 12696 10642 0 _107_
rlabel metal1 4278 12342 4278 12342 0 _108_
rlabel metal1 8418 8942 8418 8942 0 _109_
rlabel metal1 8970 7344 8970 7344 0 _110_
rlabel metal1 9062 9010 9062 9010 0 _111_
rlabel metal1 9476 6290 9476 6290 0 _112_
rlabel metal2 9706 6426 9706 6426 0 _113_
rlabel metal2 10166 6460 10166 6460 0 _114_
rlabel metal1 9246 8942 9246 8942 0 _115_
rlabel metal1 9844 9146 9844 9146 0 _116_
rlabel metal1 9752 9622 9752 9622 0 _117_
rlabel metal2 9982 10030 9982 10030 0 _118_
rlabel metal2 9522 9826 9522 9826 0 _119_
rlabel metal2 8786 9316 8786 9316 0 _120_
rlabel metal1 8878 9690 8878 9690 0 _121_
rlabel metal1 9062 9520 9062 9520 0 _122_
rlabel metal1 9384 9690 9384 9690 0 _123_
rlabel metal1 9614 6834 9614 6834 0 _124_
rlabel metal1 9614 6222 9614 6222 0 _125_
rlabel metal1 9338 6222 9338 6222 0 _126_
rlabel metal2 8970 7514 8970 7514 0 _127_
rlabel metal1 9246 6902 9246 6902 0 _128_
rlabel metal1 6624 12818 6624 12818 0 _129_
rlabel metal1 6440 12750 6440 12750 0 _130_
rlabel metal1 6670 12920 6670 12920 0 _131_
rlabel metal1 6026 12682 6026 12682 0 _132_
rlabel metal1 7176 11866 7176 11866 0 _133_
rlabel metal1 7188 11662 7188 11662 0 _134_
rlabel metal2 9246 10948 9246 10948 0 _135_
rlabel metal2 10350 9724 10350 9724 0 _136_
rlabel metal1 6670 4012 6670 4012 0 _137_
rlabel metal1 8556 3978 8556 3978 0 _138_
rlabel metal1 9798 6358 9798 6358 0 _139_
rlabel metal2 2622 11968 2622 11968 0 clk_div_bypass_en_q
rlabel metal1 6670 13702 6670 13702 0 clk_gate_state_q\[0\]
rlabel metal1 6394 13974 6394 13974 0 clk_gate_state_q\[1\]
rlabel metal3 751 12988 751 12988 0 clk_i
rlabel metal1 9798 14586 9798 14586 0 clk_o
rlabel metal2 7130 1520 7130 1520 0 cycl_count_o[0]
rlabel metal2 7774 1520 7774 1520 0 cycl_count_o[1]
rlabel metal2 8418 1520 8418 1520 0 cycl_count_o[2]
rlabel metal2 13386 4913 13386 4913 0 cycl_count_o[3]
rlabel metal2 13018 7633 13018 7633 0 cycl_count_o[4]
rlabel metal2 13386 8143 13386 8143 0 cycl_count_o[5]
rlabel metal2 13386 8857 13386 8857 0 cycl_count_o[6]
rlabel metal2 13386 9503 13386 9503 0 cycl_count_o[7]
rlabel metal3 820 11628 820 11628 0 div_i[0]
rlabel metal3 751 5508 751 5508 0 div_i[1]
rlabel metal3 751 4828 751 4828 0 div_i[2]
rlabel metal3 751 6188 751 6188 0 div_i[3]
rlabel metal3 751 8908 751 8908 0 div_i[4]
rlabel metal1 1196 6290 1196 6290 0 div_i[5]
rlabel metal3 751 6868 751 6868 0 div_i[6]
rlabel metal3 1050 8228 1050 8228 0 div_i[7]
rlabel metal1 4094 13328 4094 13328 0 div_q\[0\]
rlabel metal1 6486 4590 6486 4590 0 div_q\[1\]
rlabel metal2 8326 5406 8326 5406 0 div_q\[2\]
rlabel metal2 2254 4964 2254 4964 0 div_q\[3\]
rlabel metal1 5014 8908 5014 8908 0 div_q\[4\]
rlabel metal1 5750 7820 5750 7820 0 div_q\[5\]
rlabel metal1 8234 8466 8234 8466 0 div_q\[6\]
rlabel metal2 7958 9248 7958 9248 0 div_q\[7\]
rlabel metal1 6302 14450 6302 14450 0 div_ready_o
rlabel metal1 6302 14382 6302 14382 0 div_valid_i
rlabel metal1 7176 14382 7176 14382 0 en_i
rlabel metal1 10304 12818 10304 12818 0 even_clk
rlabel metal1 6108 13498 6108 13498 0 gate_en_d
rlabel metal1 8050 13328 8050 13328 0 gate_en_q
rlabel metal2 7038 13702 7038 13702 0 gate_is_open_q
rlabel metal1 9844 12682 9844 12682 0 i_clk_gate.clk_en
rlabel metal1 8418 13328 8418 13328 0 i_clk_gate.en_i
rlabel metal1 5060 12886 5060 12886 0 i_clk_mux.clk_sel_i
rlabel metal2 9522 12036 9522 12036 0 i_odd_clk_xor.clk1_i
rlabel metal1 1702 11764 1702 11764 0 net1
rlabel metal1 6440 14246 6440 14246 0 net10
rlabel metal1 7636 14246 7636 14246 0 net11
rlabel metal2 13294 3774 13294 3774 0 net12
rlabel metal1 8648 13294 8648 13294 0 net13
rlabel metal2 10350 14212 10350 14212 0 net14
rlabel metal2 10074 5406 10074 5406 0 net15
rlabel metal1 8004 2414 8004 2414 0 net16
rlabel metal1 8786 2448 8786 2448 0 net17
rlabel metal2 13478 5406 13478 5406 0 net18
rlabel metal1 12742 6800 12742 6800 0 net19
rlabel metal1 2116 11118 2116 11118 0 net2
rlabel metal1 13064 7854 13064 7854 0 net20
rlabel metal1 13294 9962 13294 9962 0 net21
rlabel metal2 13202 10132 13202 10132 0 net22
rlabel metal1 6072 12954 6072 12954 0 net23
rlabel metal1 2438 5100 2438 5100 0 net24
rlabel metal2 2622 8806 2622 8806 0 net25
rlabel metal2 8234 7820 8234 7820 0 net26
rlabel metal2 3082 5542 3082 5542 0 net27
rlabel metal1 5474 6290 5474 6290 0 net28
rlabel metal1 7636 2414 7636 2414 0 net29
rlabel metal2 2070 5780 2070 5780 0 net3
rlabel metal1 6999 3434 6999 3434 0 net30
rlabel metal1 10265 13226 10265 13226 0 net31
rlabel metal2 12834 5508 12834 5508 0 net32
rlabel metal2 2438 3298 2438 3298 0 net33
rlabel metal1 2622 12920 2622 12920 0 net34
rlabel metal1 11546 7310 11546 7310 0 net35
rlabel metal1 2484 7378 2484 7378 0 net36
rlabel metal2 1886 7548 1886 7548 0 net37
rlabel metal2 3358 7242 3358 7242 0 net38
rlabel metal2 2530 5338 2530 5338 0 net4
rlabel metal1 2024 5678 2024 5678 0 net5
rlabel metal2 2484 7378 2484 7378 0 net6
rlabel metal1 2438 6392 2438 6392 0 net7
rlabel metal2 2622 7684 2622 7684 0 net8
rlabel metal2 2438 8670 2438 8670 0 net9
rlabel metal2 13478 4369 13478 4369 0 rst_ni
rlabel metal1 8464 14382 8464 14382 0 test_mode_en_i
<< properties >>
string FIXED_BBOX 0 0 14989 17133
<< end >>
