* NGSPICE file created from freq_psc.ext - technology: sky130A
.subckt freq_psc_16_bit VGND VPWR clk out psc[0] psc[1] psc[2] psc[3] psc[4] psc[5] psc[6] psc[7] psc[8] psc[9]
+psc[10] psc[11] psc[12] psc[13] psc[14] psc[15] rst

X_294_ counter\[14\] _104_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__and2_1
XFILLER_13_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrebuffer7 net28 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_363_ clknet_1_0__leaf_clk _001_ _028_ VGND VGND VPWR VPWR counter\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_12_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_346_ net21 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__inv_2
X_277_ counter\[8\] _092_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__or2_1
X_200_ net15 net16 net2 VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__or3_1
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_329_ net6 _157_ _110_ _111_ _112_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__o311a_1
XFILLER_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_293_ _104_ _105_ net26 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and3b_1
X_362_ clknet_1_0__leaf_clk _015_ _027_ VGND VGND VPWR VPWR counter\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_12_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_276_ counter\[7\] counter\[8\] _090_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__and3_1
X_345_ net21 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ counter\[0\] net27 counter\[2\] VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__a21o_1
X_328_ _136_ _137_ _114_ VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_5_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_16_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_292_ counter\[13\] _102_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__or2_1
XFILLER_9_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_361_ clknet_1_0__leaf_clk _014_ _026_ VGND VGND VPWR VPWR counter\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_19_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_275_ _092_ _093_ net19 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__and3b_1
X_344_ net21 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_4_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_189_ counter\[12\] VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__inv_2
X_258_ counter\[0\] counter\[1\] counter\[2\] VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__and3_1
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_327_ _115_ _116_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__nor2_1
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_291_ counter\[13\] counter\[12\] _100_ VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__and3_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_360_ clknet_1_0__leaf_clk _013_ _025_ VGND VGND VPWR VPWR counter\[7\] sky130_fd_sc_hd__dfrtp_2
XFILLER_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_274_ counter\[7\] _090_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__or2_1
X_343_ net21 VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_20_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_188_ counter\[13\] VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__inv_2
X_257_ _049_ net20 _081_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__and3_1
X_326_ _118_ _135_ _115_ _117_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__o211a_1
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_309_ _147_ net15 net16 _152_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__o22ai_1
XFILLER_1_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ _102_ _103_ net19 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and3b_1
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_273_ counter\[7\] _090_ VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__and2_1
X_342_ net22 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_187_ net7 VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__inv_2
XFILLER_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_256_ counter\[0\] net28 VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__or2_1
X_325_ _120_ _134_ _119_ VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__a21oi_1
Xclkload0 clknet_1_0__leaf_clk VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__clkinv_2
X_308_ counter\[9\] _153_ _152_ net16 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__a2bb2o_1
X_239_ counter\[15\] _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nand2_1
XFILLER_20_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_341_ net22 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
X_272_ _090_ _091_ net20 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and3b_1
XFILLER_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_324_ _122_ _133_ _121_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_186_ net4 VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__inv_2
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_255_ _145_ net26 VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and2_4
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_238_ net7 _063_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__xnor2_1
X_307_ counter\[9\] _153_ _154_ counter\[10\] _116_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__a221oi_2
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_340_ net22 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__inv_2
X_271_ counter\[6\] _088_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__or2_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_185_ net3 VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__inv_2
X_323_ _124_ _130_ _132_ _123_ VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__a31o_1
X_254_ _076_ _075_ _079_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__o21a_4
XFILLER_2_105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_237_ net6 net25 VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__nor2_1
X_306_ counter\[11\] _155_ VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__and2_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_11_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_270_ counter\[6\] counter\[4\] counter\[5\] _084_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__and4_1
XFILLER_4_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_322_ _127_ _128_ _131_ _125_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__o211ai_1
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_184_ net2 VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__inv_2
X_253_ _065_ _067_ _078_ _069_ VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a31o_1
X_236_ _059_ counter\[13\] _060_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__and3_1
X_305_ _154_ counter\[10\] _155_ counter\[11\] VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__o22a_1
XFILLER_1_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ net10 _044_ _160_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a21boi_1
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_13_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_183_ counter\[8\] VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__inv_2
X_252_ _061_ _068_ _077_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__or3_1
X_321_ _126_ _129_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__nor2_1
X_235_ _059_ _060_ counter\[13\] VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a21oi_1
X_304_ _111_ _113_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__nand2b_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_218_ net1 net8 net9 VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__or3_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_182_ net14 VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__inv_2
X_251_ counter\[12\] _056_ _062_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__a21oi_1
X_320_ _125_ _126_ VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__nand2_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_234_ net4 _172_ net5 VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__o21ai_1
X_303_ net6 _157_ _158_ net5 _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__o221a_1
X_217_ counter\[5\] _039_ _042_ counter\[4\] VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__a22o_1
Xoutput18 net18 VGND VGND VPWR VPWR out sky130_fd_sc_hd__buf_2
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_15_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_181_ net13 VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_18_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout20 _080_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_6
X_250_ _068_ _070_ _069_ _065_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__or4b_4
XTAP_TAPCELL_ROW_0_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_302_ _156_ counter\[14\] counter\[15\] VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__a21oi_1
X_233_ _172_ net4 net5 VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__or3_4
XTAP_TAPCELL_ROW_19_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_216_ _161_ _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__and2b_1
XFILLER_18_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ net11 VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__inv_2
Xfanout21 net17 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
XFILLER_13_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_232_ counter\[12\] _056_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__and2_1
X_301_ net6 _157_ _158_ net5 _110_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__a221o_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_215_ net11 _160_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nand2_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout22 net17 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_0_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_300_ _156_ counter\[14\] VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__nor2_1
X_231_ counter\[12\] _056_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nor2_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput1 psc[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_214_ counter\[6\] _036_ _039_ counter\[5\] VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__o22a_1
XFILLER_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_230_ _155_ net23 VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__xnor2_1
X_359_ clknet_1_1__leaf_clk _012_ _024_ VGND VGND VPWR VPWR counter\[6\] sky130_fd_sc_hd__dfrtp_1
Xinput2 psc[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_7_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_213_ net12 _161_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_21_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_358_ clknet_1_1__leaf_clk _011_ _023_ VGND VGND VPWR VPWR counter\[5\] sky130_fd_sc_hd__dfrtp_2
Xinput3 psc[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ counter\[12\] _100_ VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__or2_1
X_212_ counter\[6\] _036_ _037_ counter\[7\] VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_6_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_357_ clknet_1_1__leaf_clk _010_ _022_ VGND VGND VPWR VPWR counter\[4\] sky130_fd_sc_hd__dfrtp_4
X_288_ counter\[12\] _100_ VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__and2_1
Xinput4 psc[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_211_ net14 _035_ _163_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21oi_1
XFILLER_19_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_6_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 psc[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_356_ clknet_1_1__leaf_clk _009_ _021_ VGND VGND VPWR VPWR counter\[3\] sky130_fd_sc_hd__dfrtp_2
X_287_ _100_ _101_ net19 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__and3b_1
XFILLER_19_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_210_ _150_ _034_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__xnor2_1
X_339_ net22 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__inv_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_355_ clknet_1_1__leaf_clk _008_ _020_ VGND VGND VPWR VPWR counter\[2\] sky130_fd_sc_hd__dfrtp_1
X_286_ counter\[9\] counter\[10\] _094_ counter\[11\] VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__a31o_1
Xinput6 psc[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_338_ net22 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__inv_2
X_269_ _088_ _089_ net20 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__and3b_1
XFILLER_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_14_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_354_ clknet_1_1__leaf_clk _007_ _019_ VGND VGND VPWR VPWR counter\[1\] sky130_fd_sc_hd__dfrtp_2
X_285_ counter\[11\] counter\[10\] _096_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__and3_1
Xinput7 psc[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_2_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_199_ counter\[9\] _165_ _166_ counter\[8\] _164_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__a32o_1
X_268_ counter\[4\] _084_ counter\[5\] VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__a21o_1
X_337_ net21 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__inv_2
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput10 psc[3] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_353_ clknet_1_1__leaf_clk _000_ _018_ VGND VGND VPWR VPWR counter\[0\] sky130_fd_sc_hd__dfrtp_2
X_284_ net26 _098_ _099_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__and3_1
Xinput8 psc[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_6
X_198_ net15 _160_ net24 net16 VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__o31ai_1
X_267_ counter\[4\] counter\[5\] _084_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__and3_1
X_336_ net21 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__inv_2
XFILLER_2_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput11 psc[4] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_6
X_319_ net10 counter\[2\] VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__and2b_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_12_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout19 _080_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_6
XFILLER_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_352_ clknet_1_1__leaf_clk _016_ _017_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
Xinput9 psc[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_283_ counter\[10\] _096_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__or2_1
XFILLER_14_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_197_ net15 net16 _160_ _162_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__or4_2
X_266_ net20 _086_ _087_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__and3_1
X_335_ _138_ _139_ _144_ _142_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__o22a_1
XFILLER_21_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 psc[5] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
X_249_ _175_ _055_ _074_ _071_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__o31a_1
X_318_ _145_ net8 _146_ net9 VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__o22a_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_351_ net22 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__inv_2
X_282_ counter\[10\] _096_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__nand2_1
X_334_ _114_ _115_ _117_ _143_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__nand4b_1
X_196_ net15 _163_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__xnor2_1
X_265_ counter\[4\] _084_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_6_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 psc[6] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_6
X_179_ net12 VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__inv_2
X_248_ _167_ _072_ _073_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__nand3b_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_317_ _146_ net9 VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__and2_1
XFILLER_17_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_350_ net22 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
X_281_ _096_ _097_ net26 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__and3b_1
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_195_ _160_ _162_ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__nor2_1
XFILLER_2_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_264_ counter\[4\] _084_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__nand2_1
X_333_ _119_ _123_ _124_ _128_ VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__and4bb_1
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput14 psc[7] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
X_247_ counter\[8\] _164_ _169_ counter\[10\] VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__o22a_1
X_316_ counter\[2\] net10 VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__and2b_1
X_178_ counter\[7\] VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__inv_2
XFILLER_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_280_ counter\[9\] _094_ VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_14_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_194_ net13 net11 net12 net14 VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__or4_4
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_263_ _084_ _085_ net20 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__and3b_1
X_332_ _126_ _141_ _129_ _125_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__or4b_4
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 psc[8] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
X_246_ counter\[11\] _174_ _037_ counter\[7\] _170_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__o221a_1
X_315_ counter\[3\] _149_ VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__nand2_1
X_177_ net28 VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__inv_2
XFILLER_7_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_229_ _040_ _054_ _038_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__a21oi_1
XFILLER_8_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_193_ net11 _160_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__nor2_1
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262_ counter\[3\] _082_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__or2_1
X_331_ _118_ _140_ _121_ _122_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__or4b_1
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput16 psc[9] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_314_ counter\[3\] _149_ counter\[4\] _148_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__o22a_1
X_245_ counter\[11\] _174_ _175_ _171_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__o22ai_1
X_176_ counter\[0\] VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__inv_2
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_228_ _046_ _053_ _043_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__a21o_1
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_192_ net8 net1 net9 net10 VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__or4_4
X_261_ counter\[0\] counter\[1\] counter\[2\] counter\[3\] VGND VGND VPWR VPWR _084_
+ sky130_fd_sc_hd__and4_1
X_330_ _145_ net8 _147_ net15 _127_ VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__a221o_1
X_313_ _148_ counter\[4\] counter\[5\] _150_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__a22o_1
Xinput17 rst VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
X_244_ _057_ _058_ _061_ _062_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__or4_4
X_227_ counter\[3\] _045_ _048_ _052_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a22o_1
XFILLER_8_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XTAP_TAPCELL_ROW_1_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _082_ _083_ net20 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__and3b_1
XFILLER_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ net1 net8 VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__or2_1
XFILLER_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_312_ _151_ counter\[6\] counter\[5\] _150_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__o22a_1
X_243_ counter\[15\] _064_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_1_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_226_ counter\[0\] net29 _159_ _050_ _051_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__a221o_1
X_209_ net13 _034_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__or2_1
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ net21 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_11_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_311_ _151_ counter\[6\] VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__and2_1
X_242_ counter\[14\] _066_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__xnor2_1
XFILLER_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_225_ counter\[2\] _044_ _047_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__and3_1
XFILLER_3_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclone4 _080_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_6
X_208_ net12 net11 _160_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__or3_1
XFILLER_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_310_ _147_ net15 VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__nand2_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_241_ counter\[14\] _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand2_1
XFILLER_11_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_224_ net1 _145_ net8 _146_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__o211ai_1
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_207_ counter\[10\] _169_ _174_ counter\[11\] VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_17_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_240_ net6 net25 VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__xor2_1
Xrebuffer1 _172_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XFILLER_11_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_223_ counter\[0\] net28 VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_206_ _172_ _173_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__and2_1
XFILLER_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_8_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_21_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrebuffer2 _162_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dlygate4sd1_1
X_299_ net26 _108_ _109_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and3_1
XFILLER_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_368_ clknet_1_1__leaf_clk _006_ _033_ VGND VGND VPWR VPWR counter\[15\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_222_ _044_ _047_ counter\[2\] VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__a21o_1
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_205_ net2 _165_ net3 VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_298_ counter\[15\] _106_ VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__or2_1
X_367_ clknet_1_1__leaf_clk _005_ _032_ VGND VGND VPWR VPWR counter\[14\] sky130_fd_sc_hd__dfrtp_2
Xrebuffer3 _059_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_221_ net1 net8 net9 VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__o21ai_1
X_204_ net3 _168_ _162_ _160_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__or4_4
XFILLER_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_297_ counter\[15\] _106_ VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__nand2_1
X_366_ clknet_1_0__leaf_clk _004_ _031_ VGND VGND VPWR VPWR counter\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_220_ counter\[4\] _042_ _045_ counter\[3\] VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__o22a_1
X_349_ net21 VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_8_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_203_ counter\[10\] _169_ _170_ _167_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_18_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_296_ _106_ _107_ net19 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__and3b_1
X_365_ clknet_1_0__leaf_clk _003_ _030_ VGND VGND VPWR VPWR counter\[12\] sky130_fd_sc_hd__dfrtp_2
Xrebuffer5 counter\[1\] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlygate4sd1_1
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ net21 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__inv_2
X_279_ counter\[9\] _094_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__and2_1
X_202_ _165_ _166_ counter\[9\] VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__a21o_1
XFILLER_18_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_12_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_295_ counter\[14\] _104_ VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__or2_1
Xrebuffer6 counter\[1\] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_6
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_364_ clknet_1_0__leaf_clk _002_ _029_ VGND VGND VPWR VPWR counter\[11\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_0_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_278_ _094_ _095_ net19 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__and3b_1
X_347_ net21 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__inv_2
XFILLER_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_201_ _153_ _165_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

