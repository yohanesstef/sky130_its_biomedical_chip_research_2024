magic
tech sky130A
magscale 1 2
timestamp 1729851530
<< error_p >>
rect -32 561 32 567
rect -32 527 -20 561
rect -32 521 32 527
rect -32 -527 32 -521
rect -32 -561 -20 -527
rect -32 -567 32 -561
<< nwell >>
rect -130 -580 130 580
<< pmos >>
rect -36 -480 36 480
<< pdiff >>
rect -94 468 -36 480
rect -94 -468 -82 468
rect -48 -468 -36 468
rect -94 -480 -36 -468
rect 36 468 94 480
rect 36 -468 48 468
rect 82 -468 94 468
rect 36 -480 94 -468
<< pdiffc >>
rect -82 -468 -48 468
rect 48 -468 82 468
<< poly >>
rect -36 561 36 577
rect -36 527 -20 561
rect 20 527 36 561
rect -36 480 36 527
rect -36 -527 36 -480
rect -36 -561 -20 -527
rect 20 -561 36 -527
rect -36 -577 36 -561
<< polycont >>
rect -20 527 20 561
rect -20 -561 20 -527
<< locali >>
rect -36 527 -20 561
rect 20 527 36 561
rect -82 468 -48 484
rect -82 -484 -48 -468
rect 48 468 82 484
rect 48 -484 82 -468
rect -36 -561 -20 -527
rect 20 -561 36 -527
<< viali >>
rect -20 527 20 561
rect -82 -468 -48 468
rect 48 -468 82 468
rect -20 -561 20 -527
<< metal1 >>
rect -32 561 32 567
rect -32 527 -20 561
rect 20 527 32 561
rect -32 521 32 527
rect -88 468 -42 480
rect -88 -468 -82 468
rect -48 -468 -42 468
rect -88 -480 -42 -468
rect 42 468 88 480
rect 42 -468 48 468
rect 82 -468 88 468
rect 42 -480 88 -468
rect -32 -527 32 -521
rect -32 -561 -20 -527
rect 20 -561 32 -527
rect -32 -567 32 -561
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.8 l 0.36 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
