magic
tech sky130A
magscale 1 2
timestamp 1730521008
<< nwell >>
rect -109 -314 109 348
<< pmos >>
rect -15 -214 15 286
<< pdiff >>
rect -73 274 -15 286
rect -73 -202 -61 274
rect -27 -202 -15 274
rect -73 -214 -15 -202
rect 15 274 73 286
rect 15 -202 27 274
rect 61 -202 73 274
rect 15 -214 73 -202
<< pdiffc >>
rect -61 -202 -27 274
rect 27 -202 61 274
<< poly >>
rect -15 286 15 312
rect -15 -245 15 -214
rect -33 -261 33 -245
rect -33 -295 -17 -261
rect 17 -295 33 -261
rect -33 -311 33 -295
<< polycont >>
rect -17 -295 17 -261
<< locali >>
rect -61 274 -27 290
rect -61 -218 -27 -202
rect 27 274 61 290
rect 27 -218 61 -202
rect -33 -295 -17 -261
rect 17 -295 33 -261
<< viali >>
rect -61 -202 -27 274
rect 27 -202 61 274
<< metal1 >>
rect -67 274 -21 286
rect -67 -202 -61 274
rect -27 -202 -21 274
rect -67 -214 -21 -202
rect 21 274 67 286
rect 21 -202 27 274
rect 61 -202 67 274
rect 21 -214 67 -202
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 0 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
