* NGSPICE file created from freq_psc.ext - technology: sky130A

.subckt freq_psc_8_bit VGND VPWR clk out psc[0] psc[1] psc[2] psc[3] psc[4] psc[5] psc[6]
+ psc[7] rst
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_131_ _024_ counter\[0\] counter\[1\] _023_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__o22a_1
XFILLER_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_114_ _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_5_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ _019_ counter\[5\] VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_12_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_113_ counter\[0\] counter\[1\] counter\[2\] counter\[3\] VGND VGND VPWR VPWR _054_
+ sky130_fd_sc_hd__and4_1
Xoutput10 net10 VGND VGND VPWR VPWR out sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_0_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_112_ _051_ _053_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__and2_1
XFILLER_3_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_111_ counter\[2\] _035_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__xnor2_1
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload0 clknet_1_1__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
X_110_ _035_ _051_ _052_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__and3_1
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_099_ net5 _028_ net6 VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__o21ai_1
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_098_ counter\[3\] _032_ _038_ _039_ _041_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__o221a_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_097_ counter\[4\] _040_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__or2_1
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_149_ clknet_1_0__leaf_clk _002_ _012_ VGND VGND VPWR VPWR counter\[2\] sky130_fd_sc_hd__dfrtp_2
X_096_ _021_ _028_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__xnor2_1
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_148_ clknet_1_0__leaf_clk _001_ _011_ VGND VGND VPWR VPWR counter\[1\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_11_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_079_ net2 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_3_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_095_ counter\[2\] _027_ _033_ _032_ counter\[3\] VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__a32o_1
X_078_ net3 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
XFILLER_10_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_147_ clknet_1_0__leaf_clk _000_ _010_ VGND VGND VPWR VPWR counter\[0\] sky130_fd_sc_hd__dfrtp_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_094_ _035_ _037_ _034_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a21oi_1
X_077_ net4 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__inv_2
X_129_ _018_ counter\[6\] VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__or2_1
X_146_ clknet_1_1__leaf_clk _008_ _009_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfrtp_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_093_ net2 _025_ _036_ _026_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a31o_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_076_ net5 VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__inv_2
Xinput1 psc[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_145_ net9 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ _051_ _064_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__and2_1
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 psc[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
X_092_ net1 counter\[0\] VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2b_1
XPHY_EDGE_ROW_3_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_075_ net6 VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__inv_2
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_144_ net9 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__inv_2
X_127_ counter\[7\] _062_ VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_6_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput3 psc[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_074_ net7 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__inv_2
X_091_ counter\[0\] counter\[1\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand2_1
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_143_ net9 VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_126_ _051_ _062_ _063_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__and3_1
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ counter\[0\] counter\[1\] VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__or2_1
Xinput4 psc[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_090_ _027_ _033_ counter\[2\] VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a21oi_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_073_ net8 VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__inv_2
X_142_ net9 VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__inv_2
XFILLER_2_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_125_ counter\[6\] _059_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__or2_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_108_ counter\[0\] _051_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_0_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput5 psc[4] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
X_141_ net9 VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__inv_2
X_124_ counter\[6\] _059_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__nand2_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_107_ counter\[7\] _031_ _049_ _050_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__o22ai_4
XTAP_TAPCELL_ROW_9_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 psc[5] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_140_ net9 VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__inv_2
X_106_ counter\[7\] _031_ _048_ counter\[6\] VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_10_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ _051_ _060_ _061_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 psc[6] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_10_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_122_ counter\[4\] _054_ counter\[5\] VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a21o_1
X_105_ _042_ _045_ _048_ counter\[6\] _046_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__o221a_1
XFILLER_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput8 psc[7] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_1_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_104_ _030_ _047_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and2b_1
X_121_ _059_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__inv_2
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput9 net11 VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_11_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_120_ counter\[5\] counter\[4\] _054_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__and3_1
X_103_ net7 _029_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__nand2_1
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 rst VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_2_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_102_ counter\[5\] _044_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__or2_1
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold2 counter\[7\] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_101_ counter\[4\] _040_ _044_ counter\[5\] VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__a22o_1
XFILLER_8_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_100_ _029_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__and2_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_9_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_089_ net1 net2 net3 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__o21ai_1
XFILLER_8_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_088_ _022_ _027_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_7_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ net8 _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__xnor2_2
X_139_ net9 VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__inv_2
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_086_ net7 _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_13_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_138_ net9 VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_1_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ net6 net5 _028_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__or3_1
X_154_ clknet_1_1__leaf_clk _007_ _017_ VGND VGND VPWR VPWR counter\[7\] sky130_fd_sc_hd__dfrtp_2
X_137_ _065_ _072_ net12 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a21oi_1
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_084_ net4 net3 net1 net2 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__or4_4
X_136_ _019_ counter\[5\] counter\[6\] _018_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__a221o_1
XFILLER_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_153_ clknet_1_1__leaf_clk _006_ _016_ VGND VGND VPWR VPWR counter\[6\] sky130_fd_sc_hd__dfrtp_1
X_119_ _051_ _057_ _058_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__and3_1
X_083_ net3 net1 net2 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__or3_1
X_152_ clknet_1_1__leaf_clk _005_ _015_ VGND VGND VPWR VPWR counter\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_135_ _020_ counter\[4\] _069_ _070_ _066_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__o221a_1
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_118_ counter\[4\] _054_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__or2_1
XFILLER_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_082_ net1 net2 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nor2_1
X_134_ _021_ counter\[3\] counter\[4\] _020_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__a22o_1
X_151_ clknet_1_0__leaf_clk _004_ _014_ VGND VGND VPWR VPWR counter\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_9_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_117_ counter\[4\] _054_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_081_ net9 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__inv_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_150_ clknet_1_0__leaf_clk _003_ _013_ VGND VGND VPWR VPWR counter\[3\] sky130_fd_sc_hd__dfrtp_1
X_133_ _022_ counter\[2\] counter\[3\] _021_ _068_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__o221a_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_116_ _051_ _055_ _056_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__and3_1
X_132_ _023_ counter\[1\] counter\[2\] _022_ _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__a221o_1
X_080_ counter\[1\] VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__inv_2
X_115_ counter\[0\] counter\[1\] counter\[2\] counter\[3\] VGND VGND VPWR VPWR _056_
+ sky130_fd_sc_hd__a31o_1
.ends

