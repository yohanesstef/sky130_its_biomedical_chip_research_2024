magic
tech sky130A
magscale 1 2
timestamp 1729681600
<< checkpaint >>
rect -3932 -3932 20538 22682
<< viali >>
rect 8493 16065 8527 16099
rect 9321 16065 9355 16099
rect 9873 16065 9907 16099
rect 10333 16065 10367 16099
rect 10609 16065 10643 16099
rect 11069 16065 11103 16099
rect 11713 16065 11747 16099
rect 10057 15997 10091 16031
rect 10149 15929 10183 15963
rect 8677 15861 8711 15895
rect 9137 15861 9171 15895
rect 9689 15861 9723 15895
rect 10425 15861 10459 15895
rect 11253 15861 11287 15895
rect 11897 15861 11931 15895
rect 8125 15589 8159 15623
rect 9229 15589 9263 15623
rect 12173 15589 12207 15623
rect 8585 15521 8619 15555
rect 10057 15521 10091 15555
rect 11069 15521 11103 15555
rect 11345 15521 11379 15555
rect 8309 15453 8343 15487
rect 8401 15453 8435 15487
rect 8677 15453 8711 15487
rect 8953 15453 8987 15487
rect 9597 15453 9631 15487
rect 9689 15453 9723 15487
rect 9965 15453 9999 15487
rect 10241 15453 10275 15487
rect 10333 15453 10367 15487
rect 11161 15453 11195 15487
rect 11253 15453 11287 15487
rect 11529 15453 11563 15487
rect 11621 15453 11655 15487
rect 9229 15385 9263 15419
rect 9321 15385 9355 15419
rect 11897 15385 11931 15419
rect 9045 15317 9079 15351
rect 9505 15317 9539 15351
rect 9873 15317 9907 15351
rect 10517 15317 10551 15351
rect 11805 15317 11839 15351
rect 12357 15317 12391 15351
rect 9873 15113 9907 15147
rect 11713 15113 11747 15147
rect 8309 15045 8343 15079
rect 8769 15045 8803 15079
rect 8953 15045 8987 15079
rect 9045 15045 9079 15079
rect 10057 15045 10091 15079
rect 12081 15045 12115 15079
rect 12173 15045 12207 15079
rect 8217 14977 8251 15011
rect 9142 14977 9176 15011
rect 9321 14977 9355 15011
rect 9414 14977 9448 15011
rect 9689 14977 9723 15011
rect 9781 14977 9815 15011
rect 11805 14977 11839 15011
rect 11897 14977 11931 15011
rect 12357 14977 12391 15011
rect 12449 14977 12483 15011
rect 12725 14977 12759 15011
rect 12909 14977 12943 15011
rect 13001 14977 13035 15011
rect 13093 14977 13127 15011
rect 13277 14977 13311 15011
rect 13369 14977 13403 15011
rect 6377 14909 6411 14943
rect 6653 14909 6687 14943
rect 8125 14909 8159 14943
rect 9045 14909 9079 14943
rect 11161 14909 11195 14943
rect 12817 14909 12851 14943
rect 10793 14841 10827 14875
rect 11529 14841 11563 14875
rect 12633 14841 12667 14875
rect 10057 14773 10091 14807
rect 10701 14773 10735 14807
rect 3985 14569 4019 14603
rect 7389 14569 7423 14603
rect 8401 14569 8435 14603
rect 11621 14569 11655 14603
rect 2237 14501 2271 14535
rect 1777 14365 1811 14399
rect 2605 14365 2639 14399
rect 7297 14365 7331 14399
rect 8309 14365 8343 14399
rect 10701 14365 10735 14399
rect 10793 14365 10827 14399
rect 10977 14365 11011 14399
rect 11069 14365 11103 14399
rect 11529 14365 11563 14399
rect 11713 14365 11747 14399
rect 3953 14297 3987 14331
rect 4169 14297 4203 14331
rect 2697 14229 2731 14263
rect 3801 14229 3835 14263
rect 10517 14229 10551 14263
rect 5717 14025 5751 14059
rect 6837 14025 6871 14059
rect 9137 14025 9171 14059
rect 14933 14025 14967 14059
rect 3801 13957 3835 13991
rect 5917 13957 5951 13991
rect 7021 13957 7055 13991
rect 7849 13957 7883 13991
rect 8093 13957 8127 13991
rect 8309 13957 8343 13991
rect 9873 13957 9907 13991
rect 14657 13957 14691 13991
rect 3249 13889 3283 13923
rect 3525 13889 3559 13923
rect 6009 13889 6043 13923
rect 6561 13889 6595 13923
rect 6745 13889 6779 13923
rect 7481 13889 7515 13923
rect 7665 13889 7699 13923
rect 8769 13889 8803 13923
rect 8953 13889 8987 13923
rect 9045 13889 9079 13923
rect 14565 13889 14599 13923
rect 14841 13889 14875 13923
rect 1501 13821 1535 13855
rect 2973 13821 3007 13855
rect 6101 13821 6135 13855
rect 9505 13821 9539 13855
rect 12725 13821 12759 13855
rect 14473 13821 14507 13855
rect 7389 13753 7423 13787
rect 7941 13753 7975 13787
rect 10057 13753 10091 13787
rect 5273 13685 5307 13719
rect 5549 13685 5583 13719
rect 5733 13685 5767 13719
rect 6377 13685 6411 13719
rect 7021 13685 7055 13719
rect 8125 13685 8159 13719
rect 8953 13685 8987 13719
rect 9873 13685 9907 13719
rect 12982 13685 13016 13719
rect 2421 13481 2455 13515
rect 3801 13481 3835 13515
rect 4629 13481 4663 13515
rect 7205 13481 7239 13515
rect 7481 13481 7515 13515
rect 12541 13481 12575 13515
rect 12909 13481 12943 13515
rect 14657 13481 14691 13515
rect 2881 13413 2915 13447
rect 7021 13413 7055 13447
rect 8125 13413 8159 13447
rect 11253 13413 11287 13447
rect 11713 13413 11747 13447
rect 12725 13413 12759 13447
rect 5273 13345 5307 13379
rect 5549 13345 5583 13379
rect 9781 13345 9815 13379
rect 1409 13277 1443 13311
rect 2237 13277 2271 13311
rect 2605 13277 2639 13311
rect 2697 13277 2731 13311
rect 2973 13277 3007 13311
rect 3985 13277 4019 13311
rect 4150 13277 4184 13311
rect 4267 13277 4301 13311
rect 4445 13277 4479 13311
rect 4537 13277 4571 13311
rect 7113 13277 7147 13311
rect 7297 13277 7331 13311
rect 7665 13277 7699 13311
rect 7757 13277 7791 13311
rect 8309 13277 8343 13311
rect 8493 13277 8527 13311
rect 9505 13277 9539 13311
rect 11529 13277 11563 13311
rect 11805 13277 11839 13311
rect 12173 13277 12207 13311
rect 12817 13277 12851 13311
rect 13001 13277 13035 13311
rect 14841 13277 14875 13311
rect 15117 13277 15151 13311
rect 8401 13209 8435 13243
rect 11437 13209 11471 13243
rect 1593 13141 1627 13175
rect 4353 13141 4387 13175
rect 8677 13141 8711 13175
rect 12541 13141 12575 13175
rect 14933 13141 14967 13175
rect 3065 12937 3099 12971
rect 7481 12937 7515 12971
rect 10885 12937 10919 12971
rect 11529 12937 11563 12971
rect 11805 12937 11839 12971
rect 1501 12869 1535 12903
rect 2053 12869 2087 12903
rect 10425 12869 10459 12903
rect 11253 12869 11287 12903
rect 12541 12869 12575 12903
rect 14197 12869 14231 12903
rect 3249 12801 3283 12835
rect 3433 12801 3467 12835
rect 10793 12801 10827 12835
rect 11069 12801 11103 12835
rect 11713 12801 11747 12835
rect 11897 12801 11931 12835
rect 12357 12801 12391 12835
rect 12817 12801 12851 12835
rect 13001 12801 13035 12835
rect 13737 12801 13771 12835
rect 13921 12801 13955 12835
rect 14381 12801 14415 12835
rect 14473 12801 14507 12835
rect 14749 12801 14783 12835
rect 14841 12801 14875 12835
rect 2605 12733 2639 12767
rect 7113 12733 7147 12767
rect 9229 12733 9263 12767
rect 9505 12733 9539 12767
rect 13829 12733 13863 12767
rect 14933 12733 14967 12767
rect 1869 12665 1903 12699
rect 2329 12665 2363 12699
rect 7665 12665 7699 12699
rect 12081 12665 12115 12699
rect 14657 12665 14691 12699
rect 1961 12597 1995 12631
rect 2513 12597 2547 12631
rect 3249 12597 3283 12631
rect 7481 12597 7515 12631
rect 7757 12597 7791 12631
rect 10241 12597 10275 12631
rect 10425 12597 10459 12631
rect 12725 12597 12759 12631
rect 12909 12597 12943 12631
rect 2605 12393 2639 12427
rect 4261 12393 4295 12427
rect 7665 12393 7699 12427
rect 9045 12393 9079 12427
rect 11621 12393 11655 12427
rect 13921 12393 13955 12427
rect 14933 12393 14967 12427
rect 1593 12325 1627 12359
rect 1961 12325 1995 12359
rect 2145 12325 2179 12359
rect 2467 12325 2501 12359
rect 2697 12257 2731 12291
rect 3893 12257 3927 12291
rect 5089 12257 5123 12291
rect 1409 12189 1443 12223
rect 3341 12189 3375 12223
rect 3433 12189 3467 12223
rect 4537 12189 4571 12223
rect 4721 12189 4755 12223
rect 4997 12189 5031 12223
rect 6929 12189 6963 12223
rect 7113 12189 7147 12223
rect 7389 12189 7423 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 9137 12189 9171 12223
rect 9505 12189 9539 12223
rect 11345 12189 11379 12223
rect 12173 12189 12207 12223
rect 14197 12189 14231 12223
rect 14381 12189 14415 12223
rect 14473 12189 14507 12223
rect 14565 12189 14599 12223
rect 14749 12189 14783 12223
rect 1685 12121 1719 12155
rect 2329 12121 2363 12155
rect 3065 12121 3099 12155
rect 4261 12121 4295 12155
rect 4905 12121 4939 12155
rect 6837 12121 6871 12155
rect 9781 12121 9815 12155
rect 11805 12121 11839 12155
rect 11989 12121 12023 12155
rect 12449 12121 12483 12155
rect 3157 12053 3191 12087
rect 4445 12053 4479 12087
rect 4537 12053 4571 12087
rect 7113 12053 7147 12087
rect 7297 12053 7331 12087
rect 2237 11849 2271 11883
rect 3985 11849 4019 11883
rect 6193 11849 6227 11883
rect 7205 11849 7239 11883
rect 9229 11849 9263 11883
rect 11253 11849 11287 11883
rect 11989 11849 12023 11883
rect 12081 11849 12115 11883
rect 12249 11849 12283 11883
rect 12751 11849 12785 11883
rect 13829 11849 13863 11883
rect 14565 11849 14599 11883
rect 1777 11781 1811 11815
rect 4153 11781 4187 11815
rect 4353 11781 4387 11815
rect 4721 11781 4755 11815
rect 9781 11781 9815 11815
rect 12423 11781 12457 11815
rect 12541 11781 12575 11815
rect 1409 11713 1443 11747
rect 2329 11713 2363 11747
rect 2513 11713 2547 11747
rect 2789 11713 2823 11747
rect 3065 11713 3099 11747
rect 4445 11713 4479 11747
rect 6561 11713 6595 11747
rect 6837 11713 6871 11747
rect 9137 11713 9171 11747
rect 11621 11713 11655 11747
rect 11805 11713 11839 11747
rect 13921 11713 13955 11747
rect 14657 11713 14691 11747
rect 14933 11713 14967 11747
rect 2605 11645 2639 11679
rect 9505 11645 9539 11679
rect 2053 11577 2087 11611
rect 2697 11577 2731 11611
rect 3525 11577 3559 11611
rect 12909 11577 12943 11611
rect 1593 11509 1627 11543
rect 2973 11509 3007 11543
rect 4169 11509 4203 11543
rect 6469 11509 6503 11543
rect 7205 11509 7239 11543
rect 7389 11509 7423 11543
rect 12265 11509 12299 11543
rect 12725 11509 12759 11543
rect 14841 11509 14875 11543
rect 3249 11305 3283 11339
rect 6837 11305 6871 11339
rect 8769 11305 8803 11339
rect 10517 11305 10551 11339
rect 13553 11305 13587 11339
rect 14933 11305 14967 11339
rect 1593 11237 1627 11271
rect 2697 11169 2731 11203
rect 2789 11169 2823 11203
rect 4169 11169 4203 11203
rect 5089 11169 5123 11203
rect 7297 11169 7331 11203
rect 1409 11101 1443 11135
rect 2973 11101 3007 11135
rect 3065 11101 3099 11135
rect 3341 11101 3375 11135
rect 3617 11101 3651 11135
rect 4077 11101 4111 11135
rect 4261 11101 4295 11135
rect 4353 11101 4387 11135
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 7021 11101 7055 11135
rect 9137 11101 9171 11135
rect 10425 11101 10459 11135
rect 11897 11101 11931 11135
rect 11989 11101 12023 11135
rect 12081 11101 12115 11135
rect 12173 11101 12207 11135
rect 14289 11101 14323 11135
rect 14841 11101 14875 11135
rect 15117 11101 15151 11135
rect 3525 11033 3559 11067
rect 4997 11033 5031 11067
rect 5365 11033 5399 11067
rect 9045 11033 9079 11067
rect 13645 11033 13679 11067
rect 14197 11033 14231 11067
rect 2237 10965 2271 10999
rect 11713 10965 11747 10999
rect 14657 10965 14691 10999
rect 1593 10761 1627 10795
rect 2605 10761 2639 10795
rect 6469 10761 6503 10795
rect 9949 10761 9983 10795
rect 10517 10761 10551 10795
rect 4261 10693 4295 10727
rect 10149 10693 10183 10727
rect 11897 10693 11931 10727
rect 14381 10693 14415 10727
rect 14473 10693 14507 10727
rect 14841 10693 14875 10727
rect 1409 10625 1443 10659
rect 2513 10625 2547 10659
rect 2697 10625 2731 10659
rect 5273 10625 5307 10659
rect 6561 10625 6595 10659
rect 7113 10625 7147 10659
rect 10425 10625 10459 10659
rect 10517 10625 10551 10659
rect 10701 10625 10735 10659
rect 11529 10625 11563 10659
rect 12173 10625 12207 10659
rect 14289 10625 14323 10659
rect 14657 10625 14691 10659
rect 14749 10625 14783 10659
rect 2789 10557 2823 10591
rect 3341 10557 3375 10591
rect 12449 10557 12483 10591
rect 13921 10557 13955 10591
rect 3433 10489 3467 10523
rect 3893 10489 3927 10523
rect 12081 10489 12115 10523
rect 3157 10421 3191 10455
rect 3249 10421 3283 10455
rect 3801 10421 3835 10455
rect 5365 10421 5399 10455
rect 7021 10421 7055 10455
rect 9781 10421 9815 10455
rect 9965 10421 9999 10455
rect 10333 10421 10367 10455
rect 11897 10421 11931 10455
rect 14105 10421 14139 10455
rect 10885 10217 10919 10251
rect 11713 10217 11747 10251
rect 13461 10217 13495 10251
rect 14565 10217 14599 10251
rect 1869 10149 1903 10183
rect 6009 10149 6043 10183
rect 12265 10149 12299 10183
rect 4261 10081 4295 10115
rect 8769 10081 8803 10115
rect 9045 10081 9079 10115
rect 9321 10081 9355 10115
rect 10793 10081 10827 10115
rect 12725 10081 12759 10115
rect 2237 10013 2271 10047
rect 6285 10013 6319 10047
rect 6469 10013 6503 10047
rect 6561 10013 6595 10047
rect 6653 10013 6687 10047
rect 7021 10013 7055 10047
rect 11069 10013 11103 10047
rect 11253 10013 11287 10047
rect 12357 10013 12391 10047
rect 12541 10013 12575 10047
rect 13645 10013 13679 10047
rect 13921 10013 13955 10047
rect 14105 10013 14139 10047
rect 14289 10013 14323 10047
rect 14381 10013 14415 10047
rect 14657 10013 14691 10047
rect 15117 10013 15151 10047
rect 1501 9945 1535 9979
rect 4537 9945 4571 9979
rect 6929 9945 6963 9979
rect 7297 9945 7331 9979
rect 11897 9945 11931 9979
rect 1961 9877 1995 9911
rect 2053 9877 2087 9911
rect 11989 9877 12023 9911
rect 12081 9877 12115 9911
rect 13829 9877 13863 9911
rect 14933 9877 14967 9911
rect 2789 9673 2823 9707
rect 4721 9673 4755 9707
rect 4813 9673 4847 9707
rect 11989 9673 12023 9707
rect 14565 9673 14599 9707
rect 4537 9605 4571 9639
rect 7389 9605 7423 9639
rect 8953 9605 8987 9639
rect 9321 9605 9355 9639
rect 10149 9605 10183 9639
rect 1501 9537 1535 9571
rect 2237 9537 2271 9571
rect 2513 9537 2547 9571
rect 3065 9537 3099 9571
rect 3157 9537 3191 9571
rect 3341 9537 3375 9571
rect 5089 9537 5123 9571
rect 5273 9537 5307 9571
rect 6469 9537 6503 9571
rect 9413 9537 9447 9571
rect 10517 9537 10551 9571
rect 10977 9537 11011 9571
rect 11161 9537 11195 9571
rect 11621 9537 11655 9571
rect 12265 9537 12299 9571
rect 12449 9537 12483 9571
rect 13185 9537 13219 9571
rect 14657 9537 14691 9571
rect 14933 9537 14967 9571
rect 1961 9469 1995 9503
rect 2329 9469 2363 9503
rect 2789 9469 2823 9503
rect 4997 9469 5031 9503
rect 5181 9469 5215 9503
rect 6745 9469 6779 9503
rect 12633 9469 12667 9503
rect 1777 9401 1811 9435
rect 4169 9401 4203 9435
rect 12173 9401 12207 9435
rect 2237 9333 2271 9367
rect 2697 9333 2731 9367
rect 2973 9333 3007 9367
rect 3157 9333 3191 9367
rect 4537 9333 4571 9367
rect 11069 9333 11103 9367
rect 11989 9333 12023 9367
rect 13277 9333 13311 9367
rect 14841 9333 14875 9367
rect 2237 9129 2271 9163
rect 2973 9129 3007 9163
rect 12081 9129 12115 9163
rect 14933 9129 14967 9163
rect 2145 9061 2179 9095
rect 2697 9061 2731 9095
rect 9045 9061 9079 9095
rect 2513 8993 2547 9027
rect 4629 8993 4663 9027
rect 6285 8993 6319 9027
rect 12173 8993 12207 9027
rect 12449 8993 12483 9027
rect 13921 8993 13955 9027
rect 1409 8925 1443 8959
rect 2329 8925 2363 8959
rect 2605 8925 2639 8959
rect 2789 8925 2823 8959
rect 4905 8925 4939 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 5825 8925 5859 8959
rect 5917 8925 5951 8959
rect 8953 8925 8987 8959
rect 9597 8925 9631 8959
rect 9781 8925 9815 8959
rect 10793 8925 10827 8959
rect 11621 8925 11655 8959
rect 11897 8925 11931 8959
rect 14289 8925 14323 8959
rect 14381 8925 14415 8959
rect 14657 8925 14691 8959
rect 15117 8901 15151 8935
rect 1777 8857 1811 8891
rect 4997 8857 5031 8891
rect 6193 8857 6227 8891
rect 6561 8857 6595 8891
rect 11345 8857 11379 8891
rect 11713 8857 11747 8891
rect 14473 8857 14507 8891
rect 1593 8789 1627 8823
rect 4813 8789 4847 8823
rect 5181 8789 5215 8823
rect 8033 8789 8067 8823
rect 14105 8789 14139 8823
rect 1777 8585 1811 8619
rect 4077 8585 4111 8619
rect 4813 8585 4847 8619
rect 4981 8585 5015 8619
rect 7113 8585 7147 8619
rect 7481 8585 7515 8619
rect 11345 8585 11379 8619
rect 11687 8585 11721 8619
rect 13829 8585 13863 8619
rect 14473 8585 14507 8619
rect 14933 8585 14967 8619
rect 2237 8517 2271 8551
rect 2881 8517 2915 8551
rect 5181 8517 5215 8551
rect 6469 8517 6503 8551
rect 8493 8517 8527 8551
rect 11897 8517 11931 8551
rect 13461 8517 13495 8551
rect 1409 8449 1443 8483
rect 5917 8449 5951 8483
rect 6377 8449 6411 8483
rect 6561 8449 6595 8483
rect 7113 8449 7147 8483
rect 7297 8449 7331 8483
rect 7573 8449 7607 8483
rect 7757 8449 7791 8483
rect 8033 8449 8067 8483
rect 13737 8449 13771 8483
rect 14013 8449 14047 8483
rect 14197 8449 14231 8483
rect 14289 8449 14323 8483
rect 14565 8449 14599 8483
rect 14841 8449 14875 8483
rect 15117 8449 15151 8483
rect 3028 8381 3062 8415
rect 3249 8381 3283 8415
rect 3617 8381 3651 8415
rect 3709 8381 3743 8415
rect 3985 8381 4019 8415
rect 4194 8381 4228 8415
rect 5641 8381 5675 8415
rect 9597 8381 9631 8415
rect 9873 8381 9907 8415
rect 1869 8313 1903 8347
rect 3157 8313 3191 8347
rect 4353 8313 4387 8347
rect 7849 8313 7883 8347
rect 11529 8313 11563 8347
rect 1593 8245 1627 8279
rect 4997 8245 5031 8279
rect 11713 8245 11747 8279
rect 14749 8245 14783 8279
rect 4169 8041 4203 8075
rect 5089 8041 5123 8075
rect 5273 8041 5307 8075
rect 5733 8041 5767 8075
rect 7665 8041 7699 8075
rect 9597 8041 9631 8075
rect 10701 8041 10735 8075
rect 11253 8041 11287 8075
rect 14657 8041 14691 8075
rect 14933 8041 14967 8075
rect 3065 7973 3099 8007
rect 4353 7973 4387 8007
rect 5365 7905 5399 7939
rect 8033 7905 8067 7939
rect 8677 7905 8711 7939
rect 14197 7905 14231 7939
rect 1409 7837 1443 7871
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 3341 7837 3375 7871
rect 3801 7837 3835 7871
rect 7849 7837 7883 7871
rect 8493 7837 8527 7871
rect 8769 7837 8803 7871
rect 8953 7837 8987 7871
rect 9873 7837 9907 7871
rect 9965 7837 9999 7871
rect 10221 7837 10255 7871
rect 10609 7837 10643 7871
rect 11069 7837 11103 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 14473 7837 14507 7871
rect 15117 7837 15151 7871
rect 4905 7769 4939 7803
rect 5105 7769 5139 7803
rect 8309 7769 8343 7803
rect 9321 7769 9355 7803
rect 9438 7769 9472 7803
rect 10057 7769 10091 7803
rect 10885 7769 10919 7803
rect 1593 7701 1627 7735
rect 1869 7701 1903 7735
rect 2145 7701 2179 7735
rect 3249 7701 3283 7735
rect 3433 7701 3467 7735
rect 3617 7701 3651 7735
rect 4169 7701 4203 7735
rect 5733 7701 5767 7735
rect 5917 7701 5951 7735
rect 9229 7701 9263 7735
rect 9689 7701 9723 7735
rect 2053 7497 2087 7531
rect 3065 7497 3099 7531
rect 3709 7497 3743 7531
rect 5733 7497 5767 7531
rect 6377 7497 6411 7531
rect 8861 7497 8895 7531
rect 9137 7497 9171 7531
rect 3801 7429 3835 7463
rect 5549 7429 5583 7463
rect 7849 7429 7883 7463
rect 8375 7429 8409 7463
rect 9321 7429 9355 7463
rect 13645 7429 13679 7463
rect 1501 7361 1535 7395
rect 1777 7361 1811 7395
rect 1869 7361 1903 7395
rect 2697 7361 2731 7395
rect 2881 7361 2915 7395
rect 3341 7361 3375 7395
rect 3525 7361 3559 7395
rect 3985 7361 4019 7395
rect 4077 7361 4111 7395
rect 5365 7361 5399 7395
rect 8493 7361 8527 7395
rect 8585 7361 8619 7395
rect 8677 7361 8711 7395
rect 9505 7361 9539 7395
rect 10333 7361 10367 7395
rect 11713 7361 11747 7395
rect 13737 7361 13771 7395
rect 14473 7361 14507 7395
rect 14749 7361 14783 7395
rect 2145 7293 2179 7327
rect 2605 7293 2639 7327
rect 8125 7293 8159 7327
rect 8217 7293 8251 7327
rect 11989 7293 12023 7327
rect 1593 7225 1627 7259
rect 2421 7225 2455 7259
rect 3801 7225 3835 7259
rect 14657 7225 14691 7259
rect 2789 7157 2823 7191
rect 3341 7157 3375 7191
rect 13461 7157 13495 7191
rect 14841 7157 14875 7191
rect 3893 6953 3927 6987
rect 5457 6953 5491 6987
rect 5733 6953 5767 6987
rect 8401 6953 8435 6987
rect 8585 6953 8619 6987
rect 11713 6953 11747 6987
rect 12081 6953 12115 6987
rect 12265 6953 12299 6987
rect 2053 6885 2087 6919
rect 8033 6885 8067 6919
rect 1777 6817 1811 6851
rect 2237 6817 2271 6851
rect 5089 6817 5123 6851
rect 6929 6817 6963 6851
rect 9321 6817 9355 6851
rect 12633 6817 12667 6851
rect 13369 6817 13403 6851
rect 3985 6749 4019 6783
rect 5273 6749 5307 6783
rect 6837 6749 6871 6783
rect 9505 6749 9539 6783
rect 12909 6749 12943 6783
rect 13001 6749 13035 6783
rect 13093 6749 13127 6783
rect 13185 6749 13219 6783
rect 13553 6749 13587 6783
rect 13921 6749 13955 6783
rect 14289 6749 14323 6783
rect 14381 6749 14415 6783
rect 14657 6749 14691 6783
rect 15117 6749 15151 6783
rect 5917 6681 5951 6715
rect 10241 6681 10275 6715
rect 14473 6681 14507 6715
rect 5549 6613 5583 6647
rect 5717 6613 5751 6647
rect 8401 6613 8435 6647
rect 9689 6613 9723 6647
rect 12265 6613 12299 6647
rect 12725 6613 12759 6647
rect 13645 6613 13679 6647
rect 13737 6613 13771 6647
rect 14105 6613 14139 6647
rect 14933 6613 14967 6647
rect 2513 6409 2547 6443
rect 3249 6409 3283 6443
rect 8217 6409 8251 6443
rect 9597 6409 9631 6443
rect 11621 6409 11655 6443
rect 13461 6409 13495 6443
rect 3985 6341 4019 6375
rect 5641 6341 5675 6375
rect 12357 6341 12391 6375
rect 14841 6341 14875 6375
rect 1409 6273 1443 6307
rect 2605 6273 2639 6307
rect 3433 6273 3467 6307
rect 3709 6273 3743 6307
rect 3893 6273 3927 6307
rect 4537 6273 4571 6307
rect 4721 6273 4755 6307
rect 4905 6273 4939 6307
rect 4997 6273 5031 6307
rect 5273 6273 5307 6307
rect 8493 6273 8527 6307
rect 9137 6273 9171 6307
rect 9321 6273 9355 6307
rect 11345 6273 11379 6307
rect 11713 6273 11747 6307
rect 12173 6273 12207 6307
rect 12449 6273 12483 6307
rect 13185 6273 13219 6307
rect 13645 6273 13679 6307
rect 13829 6273 13863 6307
rect 13921 6273 13955 6307
rect 14013 6273 14047 6307
rect 14197 6273 14231 6307
rect 14289 6273 14323 6307
rect 14565 6273 14599 6307
rect 14933 6273 14967 6307
rect 2053 6205 2087 6239
rect 7849 6205 7883 6239
rect 8125 6205 8159 6239
rect 8401 6205 8435 6239
rect 8769 6205 8803 6239
rect 8861 6205 8895 6239
rect 11069 6205 11103 6239
rect 1593 6137 1627 6171
rect 2329 6137 2363 6171
rect 2881 6137 2915 6171
rect 4261 6137 4295 6171
rect 4445 6137 4479 6171
rect 5825 6137 5859 6171
rect 13369 6137 13403 6171
rect 3065 6069 3099 6103
rect 5641 6069 5675 6103
rect 6377 6069 6411 6103
rect 9505 6069 9539 6103
rect 12265 6069 12299 6103
rect 14473 6069 14507 6103
rect 3801 5865 3835 5899
rect 4169 5865 4203 5899
rect 5365 5865 5399 5899
rect 8953 5865 8987 5899
rect 9965 5865 9999 5899
rect 10149 5865 10183 5899
rect 11897 5865 11931 5899
rect 14105 5865 14139 5899
rect 14841 5865 14875 5899
rect 4261 5797 4295 5831
rect 9597 5797 9631 5831
rect 13921 5797 13955 5831
rect 4077 5729 4111 5763
rect 5549 5729 5583 5763
rect 5641 5729 5675 5763
rect 12173 5729 12207 5763
rect 4537 5661 4571 5695
rect 5733 5661 5767 5695
rect 5825 5661 5859 5695
rect 6469 5661 6503 5695
rect 6837 5661 6871 5695
rect 8585 5661 8619 5695
rect 10241 5661 10275 5695
rect 14289 5661 14323 5695
rect 14381 5661 14415 5695
rect 14565 5661 14599 5695
rect 14657 5661 14691 5695
rect 14749 5661 14783 5695
rect 9137 5593 9171 5627
rect 9321 5593 9355 5627
rect 9965 5593 9999 5627
rect 10425 5593 10459 5627
rect 11713 5593 11747 5627
rect 11929 5593 11963 5627
rect 12449 5593 12483 5627
rect 4445 5525 4479 5559
rect 10609 5525 10643 5559
rect 12081 5525 12115 5559
rect 6929 5321 6963 5355
rect 8033 5321 8067 5355
rect 8861 5321 8895 5355
rect 9295 5321 9329 5355
rect 11345 5321 11379 5355
rect 12173 5321 12207 5355
rect 12541 5321 12575 5355
rect 13829 5321 13863 5355
rect 14841 5321 14875 5355
rect 8677 5253 8711 5287
rect 9505 5253 9539 5287
rect 11621 5253 11655 5287
rect 6837 5185 6871 5219
rect 7849 5185 7883 5219
rect 8033 5185 8067 5219
rect 8217 5185 8251 5219
rect 8309 5185 8343 5219
rect 8493 5185 8527 5219
rect 8769 5185 8803 5219
rect 9597 5185 9631 5219
rect 11713 5185 11747 5219
rect 12357 5185 12391 5219
rect 12633 5185 12667 5219
rect 13369 5185 13403 5219
rect 13737 5185 13771 5219
rect 14473 5185 14507 5219
rect 14749 5185 14783 5219
rect 9873 5117 9907 5151
rect 13553 5049 13587 5083
rect 14657 5049 14691 5083
rect 9045 4981 9079 5015
rect 9137 4981 9171 5015
rect 9321 4981 9355 5015
rect 3893 4777 3927 4811
rect 4537 4777 4571 4811
rect 5273 4777 5307 4811
rect 5917 4777 5951 4811
rect 7941 4777 7975 4811
rect 9965 4777 9999 4811
rect 4629 4709 4663 4743
rect 5089 4709 5123 4743
rect 10149 4709 10183 4743
rect 3341 4641 3375 4675
rect 4353 4641 4387 4675
rect 4997 4641 5031 4675
rect 1593 4573 1627 4607
rect 3617 4573 3651 4607
rect 4077 4573 4111 4607
rect 4169 4573 4203 4607
rect 4445 4573 4479 4607
rect 5549 4573 5583 4607
rect 6193 4573 6227 4607
rect 8125 4573 8159 4607
rect 8309 4573 8343 4607
rect 8401 4573 8435 4607
rect 8493 4573 8527 4607
rect 8953 4573 8987 4607
rect 9130 4573 9164 4607
rect 9597 4573 9631 4607
rect 12633 4573 12667 4607
rect 14197 4573 14231 4607
rect 1869 4505 1903 4539
rect 3525 4505 3559 4539
rect 5457 4505 5491 4539
rect 6469 4505 6503 4539
rect 9045 4505 9079 4539
rect 9965 4505 9999 4539
rect 12449 4505 12483 4539
rect 14473 4505 14507 4539
rect 5257 4437 5291 4471
rect 5917 4437 5951 4471
rect 6101 4437 6135 4471
rect 8769 4437 8803 4471
rect 12817 4437 12851 4471
rect 2789 4233 2823 4267
rect 2957 4233 2991 4267
rect 5365 4233 5399 4267
rect 5641 4233 5675 4267
rect 7573 4233 7607 4267
rect 12449 4233 12483 4267
rect 12741 4233 12775 4267
rect 3157 4165 3191 4199
rect 4629 4165 4663 4199
rect 4829 4165 4863 4199
rect 6377 4165 6411 4199
rect 6561 4165 6595 4199
rect 8769 4165 8803 4199
rect 12541 4165 12575 4199
rect 3525 4097 3559 4131
rect 3709 4097 3743 4131
rect 3801 4097 3835 4131
rect 4261 4097 4295 4131
rect 4353 4097 4387 4131
rect 5273 4097 5307 4131
rect 5457 4097 5491 4131
rect 5825 4097 5859 4131
rect 5917 4097 5951 4131
rect 7205 4097 7239 4131
rect 7297 4097 7331 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 10425 4097 10459 4131
rect 10517 4097 10551 4131
rect 12265 4097 12299 4131
rect 12449 4097 12483 4131
rect 13001 4097 13035 4131
rect 14933 4097 14967 4131
rect 15025 4097 15059 4131
rect 8493 4029 8527 4063
rect 13277 4029 13311 4063
rect 14749 4029 14783 4063
rect 4997 3961 5031 3995
rect 12909 3961 12943 3995
rect 2973 3893 3007 3927
rect 3341 3893 3375 3927
rect 4813 3893 4847 3927
rect 6745 3893 6779 3927
rect 10241 3893 10275 3927
rect 12725 3893 12759 3927
rect 5733 3689 5767 3723
rect 14933 3689 14967 3723
rect 5365 3621 5399 3655
rect 12541 3621 12575 3655
rect 4629 3553 4663 3587
rect 4077 3485 4111 3519
rect 4169 3485 4203 3519
rect 4261 3485 4295 3519
rect 4445 3485 4479 3519
rect 4537 3485 4571 3519
rect 4721 3485 4755 3519
rect 15117 3485 15151 3519
rect 5733 3417 5767 3451
rect 12265 3417 12299 3451
rect 3801 3349 3835 3383
rect 5917 3349 5951 3383
rect 12725 3349 12759 3383
rect 8493 3145 8527 3179
rect 14289 3145 14323 3179
rect 4077 3077 4111 3111
rect 5733 3077 5767 3111
rect 7849 3077 7883 3111
rect 14565 3077 14599 3111
rect 1961 3009 1995 3043
rect 3801 3009 3835 3043
rect 5825 3009 5859 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 12541 3009 12575 3043
rect 14657 3009 14691 3043
rect 2237 2941 2271 2975
rect 5549 2941 5583 2975
rect 6377 2941 6411 2975
rect 12817 2941 12851 2975
rect 3709 2805 3743 2839
rect 2053 2601 2087 2635
rect 3157 2601 3191 2635
rect 4997 2601 5031 2635
rect 6745 2601 6779 2635
rect 6929 2601 6963 2635
rect 8033 2601 8067 2635
rect 8493 2601 8527 2635
rect 7205 2533 7239 2567
rect 2237 2465 2271 2499
rect 3801 2465 3835 2499
rect 4445 2465 4479 2499
rect 2329 2397 2363 2431
rect 3249 2397 3283 2431
rect 4537 2397 4571 2431
rect 5089 2397 5123 2431
rect 6653 2397 6687 2431
rect 7113 2397 7147 2431
rect 7389 2397 7423 2431
rect 7849 2397 7883 2431
rect 8677 2397 8711 2431
rect 4721 2261 4755 2295
<< metal1 >>
rect 1104 16346 15456 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 15456 16346
rect 1104 16272 15456 16294
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 9732 16136 10364 16164
rect 9732 16124 9738 16136
rect 8386 16056 8392 16108
rect 8444 16096 8450 16108
rect 8481 16099 8539 16105
rect 8481 16096 8493 16099
rect 8444 16068 8493 16096
rect 8444 16056 8450 16068
rect 8481 16065 8493 16068
rect 8527 16065 8539 16099
rect 8481 16059 8539 16065
rect 9030 16056 9036 16108
rect 9088 16096 9094 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 9088 16068 9321 16096
rect 9088 16056 9094 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 9309 16059 9367 16065
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10336 16105 10364 16136
rect 9861 16099 9919 16105
rect 9861 16096 9873 16099
rect 9824 16068 9873 16096
rect 9824 16056 9830 16068
rect 9861 16065 9873 16068
rect 9907 16065 9919 16099
rect 9861 16059 9919 16065
rect 10321 16099 10379 16105
rect 10321 16065 10333 16099
rect 10367 16065 10379 16099
rect 10321 16059 10379 16065
rect 10410 16056 10416 16108
rect 10468 16096 10474 16108
rect 10597 16099 10655 16105
rect 10597 16096 10609 16099
rect 10468 16068 10609 16096
rect 10468 16056 10474 16068
rect 10597 16065 10609 16068
rect 10643 16065 10655 16099
rect 10597 16059 10655 16065
rect 10962 16056 10968 16108
rect 11020 16096 11026 16108
rect 11057 16099 11115 16105
rect 11057 16096 11069 16099
rect 11020 16068 11069 16096
rect 11020 16056 11026 16068
rect 11057 16065 11069 16068
rect 11103 16065 11115 16099
rect 11057 16059 11115 16065
rect 11606 16056 11612 16108
rect 11664 16096 11670 16108
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11664 16068 11713 16096
rect 11664 16056 11670 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 10045 16031 10103 16037
rect 10045 15997 10057 16031
rect 10091 15997 10103 16031
rect 10045 15991 10103 15997
rect 9950 15920 9956 15972
rect 10008 15960 10014 15972
rect 10060 15960 10088 15991
rect 10137 15963 10195 15969
rect 10137 15960 10149 15963
rect 10008 15932 10149 15960
rect 10008 15920 10014 15932
rect 10137 15929 10149 15932
rect 10183 15929 10195 15963
rect 10137 15923 10195 15929
rect 8386 15852 8392 15904
rect 8444 15892 8450 15904
rect 8665 15895 8723 15901
rect 8665 15892 8677 15895
rect 8444 15864 8677 15892
rect 8444 15852 8450 15864
rect 8665 15861 8677 15864
rect 8711 15861 8723 15895
rect 8665 15855 8723 15861
rect 8754 15852 8760 15904
rect 8812 15892 8818 15904
rect 9125 15895 9183 15901
rect 9125 15892 9137 15895
rect 8812 15864 9137 15892
rect 8812 15852 8818 15864
rect 9125 15861 9137 15864
rect 9171 15861 9183 15895
rect 9125 15855 9183 15861
rect 9214 15852 9220 15904
rect 9272 15892 9278 15904
rect 9677 15895 9735 15901
rect 9677 15892 9689 15895
rect 9272 15864 9689 15892
rect 9272 15852 9278 15864
rect 9677 15861 9689 15864
rect 9723 15892 9735 15895
rect 10042 15892 10048 15904
rect 9723 15864 10048 15892
rect 9723 15861 9735 15864
rect 9677 15855 9735 15861
rect 10042 15852 10048 15864
rect 10100 15852 10106 15904
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 10376 15864 10425 15892
rect 10376 15852 10382 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 11241 15895 11299 15901
rect 11241 15861 11253 15895
rect 11287 15892 11299 15895
rect 11606 15892 11612 15904
rect 11287 15864 11612 15892
rect 11287 15861 11299 15864
rect 11241 15855 11299 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 11882 15852 11888 15904
rect 11940 15852 11946 15904
rect 1104 15802 15456 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 15456 15802
rect 1104 15728 15456 15750
rect 8113 15623 8171 15629
rect 8113 15589 8125 15623
rect 8159 15620 8171 15623
rect 9217 15623 9275 15629
rect 8159 15592 9076 15620
rect 8159 15589 8171 15592
rect 8113 15583 8171 15589
rect 8570 15512 8576 15564
rect 8628 15512 8634 15564
rect 8294 15444 8300 15496
rect 8352 15444 8358 15496
rect 8386 15444 8392 15496
rect 8444 15444 8450 15496
rect 8665 15487 8723 15493
rect 8665 15453 8677 15487
rect 8711 15484 8723 15487
rect 8754 15484 8760 15496
rect 8711 15456 8760 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 8754 15444 8760 15456
rect 8812 15444 8818 15496
rect 8941 15487 8999 15493
rect 8941 15453 8953 15487
rect 8987 15453 8999 15487
rect 9048 15484 9076 15592
rect 9217 15589 9229 15623
rect 9263 15620 9275 15623
rect 12161 15623 12219 15629
rect 9263 15592 9720 15620
rect 9263 15589 9275 15592
rect 9217 15583 9275 15589
rect 9306 15512 9312 15564
rect 9364 15512 9370 15564
rect 9324 15484 9352 15512
rect 9692 15493 9720 15592
rect 12161 15589 12173 15623
rect 12207 15589 12219 15623
rect 12161 15583 12219 15589
rect 9766 15512 9772 15564
rect 9824 15552 9830 15564
rect 10045 15555 10103 15561
rect 10045 15552 10057 15555
rect 9824 15524 10057 15552
rect 9824 15512 9830 15524
rect 10045 15521 10057 15524
rect 10091 15521 10103 15555
rect 10045 15515 10103 15521
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11333 15555 11391 15561
rect 11333 15552 11345 15555
rect 11103 15524 11345 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 11333 15521 11345 15524
rect 11379 15521 11391 15555
rect 11882 15552 11888 15564
rect 11333 15515 11391 15521
rect 11440 15524 11888 15552
rect 9585 15487 9643 15493
rect 9585 15484 9597 15487
rect 9048 15456 9597 15484
rect 8941 15447 8999 15453
rect 9585 15453 9597 15456
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 8404 15416 8432 15444
rect 8956 15416 8984 15447
rect 9950 15444 9956 15496
rect 10008 15444 10014 15496
rect 10226 15444 10232 15496
rect 10284 15444 10290 15496
rect 10318 15444 10324 15496
rect 10376 15444 10382 15496
rect 11149 15487 11207 15493
rect 11149 15453 11161 15487
rect 11195 15453 11207 15487
rect 11149 15447 11207 15453
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15484 11299 15487
rect 11440 15484 11468 15524
rect 11882 15512 11888 15524
rect 11940 15552 11946 15564
rect 12176 15552 12204 15583
rect 11940 15524 12204 15552
rect 11940 15512 11946 15524
rect 11287 15456 11468 15484
rect 11287 15453 11299 15456
rect 11241 15447 11299 15453
rect 8404 15388 8984 15416
rect 9214 15376 9220 15428
rect 9272 15376 9278 15428
rect 9309 15419 9367 15425
rect 9309 15385 9321 15419
rect 9355 15416 9367 15419
rect 11164 15416 11192 15447
rect 11514 15444 11520 15496
rect 11572 15444 11578 15496
rect 11606 15444 11612 15496
rect 11664 15484 11670 15496
rect 12986 15484 12992 15496
rect 11664 15456 12992 15484
rect 11664 15444 11670 15456
rect 12986 15444 12992 15456
rect 13044 15444 13050 15496
rect 11330 15416 11336 15428
rect 9355 15388 10548 15416
rect 11164 15388 11336 15416
rect 9355 15385 9367 15388
rect 9309 15379 9367 15385
rect 10520 15360 10548 15388
rect 11330 15376 11336 15388
rect 11388 15416 11394 15428
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 11388 15388 11897 15416
rect 11388 15376 11394 15388
rect 11885 15385 11897 15388
rect 11931 15385 11943 15419
rect 11885 15379 11943 15385
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 9033 15351 9091 15357
rect 9033 15348 9045 15351
rect 8352 15320 9045 15348
rect 8352 15308 8358 15320
rect 9033 15317 9045 15320
rect 9079 15317 9091 15351
rect 9033 15311 9091 15317
rect 9490 15308 9496 15360
rect 9548 15308 9554 15360
rect 9858 15308 9864 15360
rect 9916 15308 9922 15360
rect 10502 15308 10508 15360
rect 10560 15308 10566 15360
rect 11790 15308 11796 15360
rect 11848 15308 11854 15360
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15348 12403 15351
rect 12710 15348 12716 15360
rect 12391 15320 12716 15348
rect 12391 15317 12403 15320
rect 12345 15311 12403 15317
rect 12710 15308 12716 15320
rect 12768 15308 12774 15360
rect 1104 15258 15456 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 15456 15258
rect 1104 15184 15456 15206
rect 9861 15147 9919 15153
rect 9861 15113 9873 15147
rect 9907 15144 9919 15147
rect 10502 15144 10508 15156
rect 9907 15116 10508 15144
rect 9907 15113 9919 15116
rect 9861 15107 9919 15113
rect 10502 15104 10508 15116
rect 10560 15104 10566 15156
rect 11701 15147 11759 15153
rect 11701 15113 11713 15147
rect 11747 15144 11759 15147
rect 11790 15144 11796 15156
rect 11747 15116 11796 15144
rect 11747 15113 11759 15116
rect 11701 15107 11759 15113
rect 11790 15104 11796 15116
rect 11848 15144 11854 15156
rect 12250 15144 12256 15156
rect 11848 15116 12256 15144
rect 11848 15104 11854 15116
rect 12250 15104 12256 15116
rect 12308 15104 12314 15156
rect 14182 15144 14188 15156
rect 12452 15116 14188 15144
rect 7282 15036 7288 15088
rect 7340 15036 7346 15088
rect 8297 15079 8355 15085
rect 8297 15045 8309 15079
rect 8343 15076 8355 15079
rect 8570 15076 8576 15088
rect 8343 15048 8576 15076
rect 8343 15045 8355 15048
rect 8297 15039 8355 15045
rect 8570 15036 8576 15048
rect 8628 15076 8634 15088
rect 8757 15079 8815 15085
rect 8757 15076 8769 15079
rect 8628 15048 8769 15076
rect 8628 15036 8634 15048
rect 8757 15045 8769 15048
rect 8803 15045 8815 15079
rect 8757 15039 8815 15045
rect 8846 15036 8852 15088
rect 8904 15076 8910 15088
rect 8941 15079 8999 15085
rect 8941 15076 8953 15079
rect 8904 15048 8953 15076
rect 8904 15036 8910 15048
rect 8941 15045 8953 15048
rect 8987 15045 8999 15079
rect 8941 15039 8999 15045
rect 9033 15079 9091 15085
rect 9033 15045 9045 15079
rect 9079 15076 9091 15079
rect 9079 15048 9996 15076
rect 9079 15045 9091 15048
rect 9033 15039 9091 15045
rect 8202 15008 8208 15020
rect 8128 14980 8208 15008
rect 5258 14900 5264 14952
rect 5316 14940 5322 14952
rect 6365 14943 6423 14949
rect 6365 14940 6377 14943
rect 5316 14912 6377 14940
rect 5316 14900 5322 14912
rect 6365 14909 6377 14912
rect 6411 14909 6423 14943
rect 6365 14903 6423 14909
rect 6638 14900 6644 14952
rect 6696 14900 6702 14952
rect 8128 14949 8156 14980
rect 8202 14968 8208 14980
rect 8260 14968 8266 15020
rect 9130 15011 9188 15017
rect 9130 15008 9142 15011
rect 8956 14980 9142 15008
rect 8113 14943 8171 14949
rect 8113 14909 8125 14943
rect 8159 14909 8171 14943
rect 8113 14903 8171 14909
rect 8956 14872 8984 14980
rect 9130 14977 9142 14980
rect 9176 14977 9188 15011
rect 9130 14971 9188 14977
rect 9306 14968 9312 15020
rect 9364 14968 9370 15020
rect 9402 15011 9460 15017
rect 9402 14977 9414 15011
rect 9448 15008 9460 15011
rect 9490 15008 9496 15020
rect 9448 14980 9496 15008
rect 9448 14977 9460 14980
rect 9402 14971 9460 14977
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 9416 14940 9444 14971
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 15008 9735 15011
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 9723 14980 9781 15008
rect 9723 14977 9735 14980
rect 9677 14971 9735 14977
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 9968 15008 9996 15048
rect 10042 15036 10048 15088
rect 10100 15036 10106 15088
rect 10686 15036 10692 15088
rect 10744 15076 10750 15088
rect 12069 15079 12127 15085
rect 12069 15076 12081 15079
rect 10744 15048 12081 15076
rect 10744 15036 10750 15048
rect 12069 15045 12081 15048
rect 12115 15045 12127 15079
rect 12069 15039 12127 15045
rect 12158 15036 12164 15088
rect 12216 15036 12222 15088
rect 10318 15008 10324 15020
rect 9968 14980 10324 15008
rect 9769 14971 9827 14977
rect 10318 14968 10324 14980
rect 10376 14968 10382 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11882 14968 11888 15020
rect 11940 14968 11946 15020
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12452 15017 12480 15116
rect 14182 15104 14188 15116
rect 14240 15104 14246 15156
rect 12728 15048 13492 15076
rect 12728 15020 12756 15048
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 12032 14980 12357 15008
rect 12032 14968 12038 14980
rect 12345 14977 12357 14980
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12437 15011 12495 15017
rect 12437 14977 12449 15011
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12710 14968 12716 15020
rect 12768 14968 12774 15020
rect 12897 15011 12955 15017
rect 12897 14977 12909 15011
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 10226 14940 10232 14952
rect 9079 14912 9444 14940
rect 9508 14912 10232 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 9508 14872 9536 14912
rect 10226 14900 10232 14912
rect 10284 14900 10290 14952
rect 11149 14943 11207 14949
rect 11149 14909 11161 14943
rect 11195 14940 11207 14943
rect 12066 14940 12072 14952
rect 11195 14912 12072 14940
rect 11195 14909 11207 14912
rect 11149 14903 11207 14909
rect 12066 14900 12072 14912
rect 12124 14900 12130 14952
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 12176 14912 12817 14940
rect 8956 14844 9536 14872
rect 9858 14832 9864 14884
rect 9916 14872 9922 14884
rect 10781 14875 10839 14881
rect 10781 14872 10793 14875
rect 9916 14844 10793 14872
rect 9916 14832 9922 14844
rect 10781 14841 10793 14844
rect 10827 14872 10839 14875
rect 11517 14875 11575 14881
rect 11517 14872 11529 14875
rect 10827 14844 11529 14872
rect 10827 14841 10839 14844
rect 10781 14835 10839 14841
rect 11517 14841 11529 14844
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 11790 14832 11796 14884
rect 11848 14872 11854 14884
rect 12176 14872 12204 14912
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 11848 14844 12204 14872
rect 11848 14832 11854 14844
rect 12250 14832 12256 14884
rect 12308 14872 12314 14884
rect 12621 14875 12679 14881
rect 12621 14872 12633 14875
rect 12308 14844 12633 14872
rect 12308 14832 12314 14844
rect 12621 14841 12633 14844
rect 12667 14841 12679 14875
rect 12621 14835 12679 14841
rect 10042 14764 10048 14816
rect 10100 14764 10106 14816
rect 10689 14807 10747 14813
rect 10689 14773 10701 14807
rect 10735 14804 10747 14807
rect 10962 14804 10968 14816
rect 10735 14776 10968 14804
rect 10735 14773 10747 14776
rect 10689 14767 10747 14773
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 12342 14764 12348 14816
rect 12400 14804 12406 14816
rect 12912 14804 12940 14971
rect 12986 14968 12992 15020
rect 13044 14968 13050 15020
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13096 14940 13124 14971
rect 13262 14968 13268 15020
rect 13320 14968 13326 15020
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15006 13415 15011
rect 13464 15006 13492 15048
rect 13403 14978 13492 15006
rect 13403 14977 13415 14978
rect 13357 14971 13415 14977
rect 14642 14940 14648 14952
rect 13096 14912 14648 14940
rect 14642 14900 14648 14912
rect 14700 14900 14706 14952
rect 12400 14776 12940 14804
rect 12400 14764 12406 14776
rect 1104 14714 15456 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 15456 14714
rect 1104 14640 15456 14662
rect 3970 14560 3976 14612
rect 4028 14560 4034 14612
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 7377 14603 7435 14609
rect 7377 14600 7389 14603
rect 7340 14572 7389 14600
rect 7340 14560 7346 14572
rect 7377 14569 7389 14572
rect 7423 14569 7435 14603
rect 7377 14563 7435 14569
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8389 14603 8447 14609
rect 8389 14600 8401 14603
rect 8352 14572 8401 14600
rect 8352 14560 8358 14572
rect 8389 14569 8401 14572
rect 8435 14569 8447 14603
rect 8389 14563 8447 14569
rect 11609 14603 11667 14609
rect 11609 14569 11621 14603
rect 11655 14600 11667 14603
rect 11974 14600 11980 14612
rect 11655 14572 11980 14600
rect 11655 14569 11667 14572
rect 11609 14563 11667 14569
rect 11974 14560 11980 14572
rect 12032 14560 12038 14612
rect 2225 14535 2283 14541
rect 2225 14501 2237 14535
rect 2271 14501 2283 14535
rect 2225 14495 2283 14501
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1728 14368 1777 14396
rect 1728 14356 1734 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 2240 14396 2268 14495
rect 11882 14492 11888 14544
rect 11940 14532 11946 14544
rect 14550 14532 14556 14544
rect 11940 14504 14556 14532
rect 11940 14492 11946 14504
rect 14550 14492 14556 14504
rect 14608 14492 14614 14544
rect 10042 14424 10048 14476
rect 10100 14464 10106 14476
rect 11790 14464 11796 14476
rect 10100 14436 11100 14464
rect 10100 14424 10106 14436
rect 2593 14399 2651 14405
rect 2593 14396 2605 14399
rect 2240 14368 2605 14396
rect 1765 14359 1823 14365
rect 2593 14365 2605 14368
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 5994 14356 6000 14408
rect 6052 14396 6058 14408
rect 7285 14399 7343 14405
rect 7285 14396 7297 14399
rect 6052 14368 7297 14396
rect 6052 14356 6058 14368
rect 7285 14365 7297 14368
rect 7331 14365 7343 14399
rect 7285 14359 7343 14365
rect 8294 14356 8300 14408
rect 8352 14356 8358 14408
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 10781 14399 10839 14405
rect 10781 14365 10793 14399
rect 10827 14365 10839 14399
rect 10781 14359 10839 14365
rect 3878 14288 3884 14340
rect 3936 14337 3942 14340
rect 3936 14331 3999 14337
rect 3936 14297 3953 14331
rect 3987 14297 3999 14331
rect 3936 14291 3999 14297
rect 4157 14331 4215 14337
rect 4157 14297 4169 14331
rect 4203 14328 4215 14331
rect 4706 14328 4712 14340
rect 4203 14300 4712 14328
rect 4203 14297 4215 14300
rect 4157 14291 4215 14297
rect 3936 14288 3942 14291
rect 4706 14288 4712 14300
rect 4764 14328 4770 14340
rect 5442 14328 5448 14340
rect 4764 14300 5448 14328
rect 4764 14288 4770 14300
rect 5442 14288 5448 14300
rect 5500 14288 5506 14340
rect 8754 14288 8760 14340
rect 8812 14328 8818 14340
rect 9766 14328 9772 14340
rect 8812 14300 9772 14328
rect 8812 14288 8818 14300
rect 9766 14288 9772 14300
rect 9824 14288 9830 14340
rect 10796 14328 10824 14359
rect 10962 14356 10968 14408
rect 11020 14356 11026 14408
rect 11072 14405 11100 14436
rect 11532 14436 11796 14464
rect 11532 14405 11560 14436
rect 11790 14424 11796 14436
rect 11848 14424 11854 14476
rect 11057 14399 11115 14405
rect 11057 14365 11069 14399
rect 11103 14365 11115 14399
rect 11057 14359 11115 14365
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14365 11575 14399
rect 11517 14359 11575 14365
rect 11698 14356 11704 14408
rect 11756 14356 11762 14408
rect 10796 14300 12434 14328
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 2685 14263 2743 14269
rect 2685 14260 2697 14263
rect 2648 14232 2697 14260
rect 2648 14220 2654 14232
rect 2685 14229 2697 14232
rect 2731 14229 2743 14263
rect 2685 14223 2743 14229
rect 3786 14220 3792 14272
rect 3844 14220 3850 14272
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 10505 14263 10563 14269
rect 10505 14260 10517 14263
rect 9732 14232 10517 14260
rect 9732 14220 9738 14232
rect 10505 14229 10517 14232
rect 10551 14229 10563 14263
rect 10505 14223 10563 14229
rect 11606 14220 11612 14272
rect 11664 14260 11670 14272
rect 12250 14260 12256 14272
rect 11664 14232 12256 14260
rect 11664 14220 11670 14232
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12406 14260 12434 14300
rect 13446 14260 13452 14272
rect 12406 14232 13452 14260
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 1104 14170 15456 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 15456 14170
rect 1104 14096 15456 14118
rect 5258 14056 5264 14068
rect 3528 14028 5264 14056
rect 2866 13988 2872 14000
rect 2530 13960 2872 13988
rect 2866 13948 2872 13960
rect 2924 13948 2930 14000
rect 3528 13929 3556 14028
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 5705 14059 5763 14065
rect 5705 14025 5717 14059
rect 5751 14056 5763 14059
rect 5751 14028 6592 14056
rect 5751 14025 5763 14028
rect 5705 14019 5763 14025
rect 3786 13948 3792 14000
rect 3844 13948 3850 14000
rect 4798 13948 4804 14000
rect 4856 13948 4862 14000
rect 5905 13991 5963 13997
rect 5905 13957 5917 13991
rect 5951 13988 5963 13991
rect 6454 13988 6460 14000
rect 5951 13960 6460 13988
rect 5951 13957 5963 13960
rect 5905 13951 5963 13957
rect 6454 13948 6460 13960
rect 6512 13948 6518 14000
rect 6564 13988 6592 14028
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6696 14028 6837 14056
rect 6696 14016 6702 14028
rect 6825 14025 6837 14028
rect 6871 14025 6883 14059
rect 6825 14019 6883 14025
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 10226 14056 10232 14068
rect 9171 14028 10232 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 6914 13988 6920 14000
rect 6564 13960 6920 13988
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7009 13991 7067 13997
rect 7009 13957 7021 13991
rect 7055 13988 7067 13991
rect 7837 13991 7895 13997
rect 7837 13988 7849 13991
rect 7055 13960 7849 13988
rect 7055 13957 7067 13960
rect 7009 13951 7067 13957
rect 7837 13957 7849 13960
rect 7883 13957 7895 13991
rect 7837 13951 7895 13957
rect 8018 13948 8024 14000
rect 8076 13997 8082 14000
rect 8076 13991 8139 13997
rect 8076 13957 8093 13991
rect 8127 13957 8139 13991
rect 8076 13951 8139 13957
rect 8076 13948 8082 13951
rect 8202 13948 8208 14000
rect 8260 13988 8266 14000
rect 8297 13991 8355 13997
rect 8297 13988 8309 13991
rect 8260 13960 8309 13988
rect 8260 13948 8266 13960
rect 8297 13957 8309 13960
rect 8343 13957 8355 13991
rect 9140 13988 9168 14019
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 13262 14016 13268 14068
rect 13320 14056 13326 14068
rect 14921 14059 14979 14065
rect 14921 14056 14933 14059
rect 13320 14028 14933 14056
rect 13320 14016 13326 14028
rect 14921 14025 14933 14028
rect 14967 14025 14979 14059
rect 14921 14019 14979 14025
rect 8297 13951 8355 13957
rect 8956 13960 9168 13988
rect 3237 13923 3295 13929
rect 3237 13889 3249 13923
rect 3283 13920 3295 13923
rect 3513 13923 3571 13929
rect 3513 13920 3525 13923
rect 3283 13892 3525 13920
rect 3283 13889 3295 13892
rect 3237 13883 3295 13889
rect 3513 13889 3525 13892
rect 3559 13889 3571 13923
rect 3513 13883 3571 13889
rect 5994 13880 6000 13932
rect 6052 13880 6058 13932
rect 6549 13923 6607 13929
rect 6549 13889 6561 13923
rect 6595 13889 6607 13923
rect 6549 13883 6607 13889
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13920 6791 13923
rect 6779 13892 7328 13920
rect 6779 13889 6791 13892
rect 6733 13883 6791 13889
rect 1489 13855 1547 13861
rect 1489 13821 1501 13855
rect 1535 13852 1547 13855
rect 1670 13852 1676 13864
rect 1535 13824 1676 13852
rect 1535 13821 1547 13824
rect 1489 13815 1547 13821
rect 1670 13812 1676 13824
rect 1728 13812 1734 13864
rect 2958 13812 2964 13864
rect 3016 13812 3022 13864
rect 6086 13812 6092 13864
rect 6144 13812 6150 13864
rect 6564 13852 6592 13883
rect 7006 13852 7012 13864
rect 6564 13824 7012 13852
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 7300 13796 7328 13892
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 7653 13923 7711 13929
rect 7653 13889 7665 13923
rect 7699 13920 7711 13923
rect 8220 13920 8248 13948
rect 7699 13892 8248 13920
rect 7699 13889 7711 13892
rect 7653 13883 7711 13889
rect 8754 13880 8760 13932
rect 8812 13880 8818 13932
rect 8956 13929 8984 13960
rect 9858 13948 9864 14000
rect 9916 13948 9922 14000
rect 14645 13991 14703 13997
rect 14645 13988 14657 13991
rect 14214 13960 14657 13988
rect 14645 13957 14657 13960
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 8941 13923 8999 13929
rect 8941 13889 8953 13923
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13889 9091 13923
rect 14553 13923 14611 13929
rect 14553 13920 14565 13923
rect 9033 13883 9091 13889
rect 14200 13892 14565 13920
rect 7558 13812 7564 13864
rect 7616 13852 7622 13864
rect 9048 13852 9076 13883
rect 7616 13824 9076 13852
rect 9493 13855 9551 13861
rect 7616 13812 7622 13824
rect 9493 13821 9505 13855
rect 9539 13852 9551 13855
rect 9539 13824 10180 13852
rect 9539 13821 9551 13824
rect 9493 13815 9551 13821
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 5500 13756 7052 13784
rect 5500 13744 5506 13756
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 5261 13719 5319 13725
rect 5261 13716 5273 13719
rect 4948 13688 5273 13716
rect 4948 13676 4954 13688
rect 5261 13685 5273 13688
rect 5307 13685 5319 13719
rect 5261 13679 5319 13685
rect 5534 13676 5540 13728
rect 5592 13676 5598 13728
rect 7024 13725 7052 13756
rect 7282 13744 7288 13796
rect 7340 13784 7346 13796
rect 7377 13787 7435 13793
rect 7377 13784 7389 13787
rect 7340 13756 7389 13784
rect 7340 13744 7346 13756
rect 7377 13753 7389 13756
rect 7423 13784 7435 13787
rect 7929 13787 7987 13793
rect 7929 13784 7941 13787
rect 7423 13756 7941 13784
rect 7423 13753 7435 13756
rect 7377 13747 7435 13753
rect 7929 13753 7941 13756
rect 7975 13753 7987 13787
rect 7929 13747 7987 13753
rect 8018 13744 8024 13796
rect 8076 13784 8082 13796
rect 9508 13784 9536 13815
rect 8076 13756 9536 13784
rect 8076 13744 8082 13756
rect 9766 13744 9772 13796
rect 9824 13784 9830 13796
rect 10045 13787 10103 13793
rect 10045 13784 10057 13787
rect 9824 13756 10057 13784
rect 9824 13744 9830 13756
rect 10045 13753 10057 13756
rect 10091 13753 10103 13787
rect 10152 13784 10180 13824
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 12713 13855 12771 13861
rect 12713 13852 12725 13855
rect 12216 13824 12725 13852
rect 12216 13812 12222 13824
rect 12713 13821 12725 13824
rect 12759 13821 12771 13855
rect 13998 13852 14004 13864
rect 12713 13815 12771 13821
rect 12820 13824 14004 13852
rect 10962 13784 10968 13796
rect 10152 13756 10968 13784
rect 10045 13747 10103 13753
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 11514 13744 11520 13796
rect 11572 13784 11578 13796
rect 12820 13784 12848 13824
rect 13998 13812 14004 13824
rect 14056 13852 14062 13864
rect 14200 13852 14228 13892
rect 14553 13889 14565 13892
rect 14599 13889 14611 13923
rect 14553 13883 14611 13889
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 14056 13824 14228 13852
rect 14461 13855 14519 13861
rect 14056 13812 14062 13824
rect 14461 13821 14473 13855
rect 14507 13852 14519 13855
rect 14844 13852 14872 13883
rect 14507 13824 14872 13852
rect 14507 13821 14519 13824
rect 14461 13815 14519 13821
rect 11572 13756 12848 13784
rect 11572 13744 11578 13756
rect 5721 13719 5779 13725
rect 5721 13685 5733 13719
rect 5767 13716 5779 13719
rect 6365 13719 6423 13725
rect 6365 13716 6377 13719
rect 5767 13688 6377 13716
rect 5767 13685 5779 13688
rect 5721 13679 5779 13685
rect 6365 13685 6377 13688
rect 6411 13685 6423 13719
rect 6365 13679 6423 13685
rect 7009 13719 7067 13725
rect 7009 13685 7021 13719
rect 7055 13716 7067 13719
rect 7098 13716 7104 13728
rect 7055 13688 7104 13716
rect 7055 13685 7067 13688
rect 7009 13679 7067 13685
rect 7098 13676 7104 13688
rect 7156 13676 7162 13728
rect 7742 13676 7748 13728
rect 7800 13716 7806 13728
rect 8113 13719 8171 13725
rect 8113 13716 8125 13719
rect 7800 13688 8125 13716
rect 7800 13676 7806 13688
rect 8113 13685 8125 13688
rect 8159 13716 8171 13719
rect 8294 13716 8300 13728
rect 8159 13688 8300 13716
rect 8159 13685 8171 13688
rect 8113 13679 8171 13685
rect 8294 13676 8300 13688
rect 8352 13676 8358 13728
rect 8938 13676 8944 13728
rect 8996 13676 9002 13728
rect 9861 13719 9919 13725
rect 9861 13685 9873 13719
rect 9907 13716 9919 13719
rect 9950 13716 9956 13728
rect 9907 13688 9956 13716
rect 9907 13685 9919 13688
rect 9861 13679 9919 13685
rect 9950 13676 9956 13688
rect 10008 13676 10014 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 12970 13719 13028 13725
rect 12970 13716 12982 13719
rect 12768 13688 12982 13716
rect 12768 13676 12774 13688
rect 12970 13685 12982 13688
rect 13016 13685 13028 13719
rect 12970 13679 13028 13685
rect 1104 13626 15456 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 15456 13626
rect 1104 13552 15456 13574
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2958 13512 2964 13524
rect 2455 13484 2964 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 3789 13515 3847 13521
rect 3789 13481 3801 13515
rect 3835 13512 3847 13515
rect 3970 13512 3976 13524
rect 3835 13484 3976 13512
rect 3835 13481 3847 13484
rect 3789 13475 3847 13481
rect 3970 13472 3976 13484
rect 4028 13472 4034 13524
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 4798 13512 4804 13524
rect 4663 13484 4804 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5994 13512 6000 13524
rect 5184 13484 6000 13512
rect 2866 13404 2872 13456
rect 2924 13404 2930 13456
rect 3050 13404 3056 13456
rect 3108 13444 3114 13456
rect 5184 13444 5212 13484
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6914 13472 6920 13524
rect 6972 13512 6978 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 6972 13484 7205 13512
rect 6972 13472 6978 13484
rect 7193 13481 7205 13484
rect 7239 13481 7251 13515
rect 7193 13475 7251 13481
rect 7466 13472 7472 13524
rect 7524 13472 7530 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 12529 13515 12587 13521
rect 10008 13484 12434 13512
rect 10008 13472 10014 13484
rect 3108 13416 5212 13444
rect 3108 13404 3114 13416
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 4890 13376 4896 13388
rect 4396 13348 4896 13376
rect 4396 13336 4402 13348
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 900 13280 1409 13308
rect 900 13268 906 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 2222 13268 2228 13320
rect 2280 13268 2286 13320
rect 2590 13268 2596 13320
rect 2648 13268 2654 13320
rect 2685 13311 2743 13317
rect 2685 13277 2697 13311
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13308 3019 13311
rect 3050 13308 3056 13320
rect 3007 13280 3056 13308
rect 3007 13277 3019 13280
rect 2961 13271 3019 13277
rect 1486 13132 1492 13184
rect 1544 13172 1550 13184
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 1544 13144 1593 13172
rect 1544 13132 1550 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 2700 13172 2728 13271
rect 3050 13268 3056 13280
rect 3108 13268 3114 13320
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 4154 13317 4160 13320
rect 4138 13311 4160 13317
rect 4138 13277 4150 13311
rect 4138 13271 4160 13277
rect 4154 13268 4160 13271
rect 4212 13268 4218 13320
rect 4246 13268 4252 13320
rect 4304 13317 4310 13320
rect 4448 13317 4476 13348
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 4304 13308 4313 13317
rect 4433 13311 4491 13317
rect 4304 13280 4349 13308
rect 4304 13271 4313 13280
rect 4433 13277 4445 13311
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 4525 13311 4583 13317
rect 4525 13277 4537 13311
rect 4571 13308 4583 13311
rect 5184 13308 5212 13416
rect 7006 13404 7012 13456
rect 7064 13444 7070 13456
rect 7558 13444 7564 13456
rect 7064 13416 7564 13444
rect 7064 13404 7070 13416
rect 5258 13336 5264 13388
rect 5316 13336 5322 13388
rect 5534 13336 5540 13388
rect 5592 13336 5598 13388
rect 7116 13317 7144 13416
rect 7558 13404 7564 13416
rect 7616 13404 7622 13456
rect 8113 13447 8171 13453
rect 8113 13413 8125 13447
rect 8159 13444 8171 13447
rect 8202 13444 8208 13456
rect 8159 13416 8208 13444
rect 8159 13413 8171 13416
rect 8113 13407 8171 13413
rect 8202 13404 8208 13416
rect 8260 13404 8266 13456
rect 11241 13447 11299 13453
rect 11241 13413 11253 13447
rect 11287 13444 11299 13447
rect 11330 13444 11336 13456
rect 11287 13416 11336 13444
rect 11287 13413 11299 13416
rect 11241 13407 11299 13413
rect 11330 13404 11336 13416
rect 11388 13404 11394 13456
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 11701 13447 11759 13453
rect 11701 13444 11713 13447
rect 11664 13416 11713 13444
rect 11664 13404 11670 13416
rect 11701 13413 11713 13416
rect 11747 13413 11759 13447
rect 11701 13407 11759 13413
rect 9766 13336 9772 13388
rect 9824 13336 9830 13388
rect 4571 13280 5212 13308
rect 7101 13311 7159 13317
rect 4571 13277 4583 13280
rect 4525 13271 4583 13277
rect 7101 13277 7113 13311
rect 7147 13277 7159 13311
rect 7101 13271 7159 13277
rect 4304 13268 4310 13271
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 2774 13200 2780 13252
rect 2832 13240 2838 13252
rect 3988 13240 4016 13268
rect 2832 13212 4016 13240
rect 2832 13200 2838 13212
rect 6086 13200 6092 13252
rect 6144 13200 6150 13252
rect 7668 13240 7696 13271
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 8297 13311 8355 13317
rect 8297 13308 8309 13311
rect 7800 13280 8309 13308
rect 7800 13268 7806 13280
rect 8297 13277 8309 13280
rect 8343 13277 8355 13311
rect 8297 13271 8355 13277
rect 8481 13311 8539 13317
rect 8481 13277 8493 13311
rect 8527 13308 8539 13311
rect 8938 13308 8944 13320
rect 8527 13280 8944 13308
rect 8527 13277 8539 13280
rect 8481 13271 8539 13277
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 11514 13268 11520 13320
rect 11572 13268 11578 13320
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13308 11851 13311
rect 11882 13308 11888 13320
rect 11839 13280 11888 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 11974 13268 11980 13320
rect 12032 13308 12038 13320
rect 12161 13311 12219 13317
rect 12161 13308 12173 13311
rect 12032 13280 12173 13308
rect 12032 13268 12038 13280
rect 12161 13277 12173 13280
rect 12207 13277 12219 13311
rect 12161 13271 12219 13277
rect 8018 13240 8024 13252
rect 7668 13212 8024 13240
rect 8018 13200 8024 13212
rect 8076 13240 8082 13252
rect 8389 13243 8447 13249
rect 8389 13240 8401 13243
rect 8076 13212 8401 13240
rect 8076 13200 8082 13212
rect 8389 13209 8401 13212
rect 8435 13209 8447 13243
rect 11425 13243 11483 13249
rect 11425 13240 11437 13243
rect 10994 13212 11437 13240
rect 8389 13203 8447 13209
rect 11425 13209 11437 13212
rect 11471 13209 11483 13243
rect 11425 13203 11483 13209
rect 3878 13172 3884 13184
rect 2700 13144 3884 13172
rect 1581 13135 1639 13141
rect 3878 13132 3884 13144
rect 3936 13172 3942 13184
rect 4341 13175 4399 13181
rect 4341 13172 4353 13175
rect 3936 13144 4353 13172
rect 3936 13132 3942 13144
rect 4341 13141 4353 13144
rect 4387 13141 4399 13175
rect 4341 13135 4399 13141
rect 8662 13132 8668 13184
rect 8720 13132 8726 13184
rect 12406 13172 12434 13484
rect 12529 13481 12541 13515
rect 12575 13512 12587 13515
rect 12897 13515 12955 13521
rect 12897 13512 12909 13515
rect 12575 13484 12909 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12897 13481 12909 13484
rect 12943 13481 12955 13515
rect 12897 13475 12955 13481
rect 14642 13472 14648 13524
rect 14700 13472 14706 13524
rect 12710 13404 12716 13456
rect 12768 13404 12774 13456
rect 12805 13311 12863 13317
rect 12805 13277 12817 13311
rect 12851 13308 12863 13311
rect 12894 13308 12900 13320
rect 12851 13280 12900 13308
rect 12851 13277 12863 13280
rect 12805 13271 12863 13277
rect 12894 13268 12900 13280
rect 12952 13268 12958 13320
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13308 13047 13311
rect 13262 13308 13268 13320
rect 13035 13280 13268 13308
rect 13035 13277 13047 13280
rect 12989 13271 13047 13277
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 14826 13268 14832 13320
rect 14884 13268 14890 13320
rect 15105 13311 15163 13317
rect 15105 13277 15117 13311
rect 15151 13308 15163 13311
rect 15194 13308 15200 13320
rect 15151 13280 15200 13308
rect 15151 13277 15163 13280
rect 15105 13271 15163 13277
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 12526 13172 12532 13184
rect 12406 13144 12532 13172
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 14918 13132 14924 13184
rect 14976 13132 14982 13184
rect 1104 13082 15456 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 15456 13082
rect 1104 13008 15456 13030
rect 3053 12971 3111 12977
rect 3053 12937 3065 12971
rect 3099 12937 3111 12971
rect 3053 12931 3111 12937
rect 7469 12971 7527 12977
rect 7469 12937 7481 12971
rect 7515 12968 7527 12971
rect 7515 12940 9812 12968
rect 7515 12937 7527 12940
rect 7469 12931 7527 12937
rect 1486 12860 1492 12912
rect 1544 12860 1550 12912
rect 1854 12860 1860 12912
rect 1912 12900 1918 12912
rect 2041 12903 2099 12909
rect 2041 12900 2053 12903
rect 1912 12872 2053 12900
rect 1912 12860 1918 12872
rect 2041 12869 2053 12872
rect 2087 12900 2099 12903
rect 2774 12900 2780 12912
rect 2087 12872 2780 12900
rect 2087 12869 2099 12872
rect 2041 12863 2099 12869
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 1504 12832 1532 12860
rect 3068 12832 3096 12931
rect 8202 12860 8208 12912
rect 8260 12860 8266 12912
rect 9784 12900 9812 12940
rect 9858 12928 9864 12980
rect 9916 12968 9922 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 9916 12940 10885 12968
rect 9916 12928 9922 12940
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 11020 12940 11529 12968
rect 11020 12928 11026 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11517 12931 11575 12937
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11793 12971 11851 12977
rect 11793 12968 11805 12971
rect 11756 12940 11805 12968
rect 11756 12928 11762 12940
rect 11793 12937 11805 12940
rect 11839 12968 11851 12971
rect 11839 12940 12204 12968
rect 11839 12937 11851 12940
rect 11793 12931 11851 12937
rect 9950 12900 9956 12912
rect 9784 12872 9956 12900
rect 9950 12860 9956 12872
rect 10008 12900 10014 12912
rect 10413 12903 10471 12909
rect 10413 12900 10425 12903
rect 10008 12872 10425 12900
rect 10008 12860 10014 12872
rect 10413 12869 10425 12872
rect 10459 12869 10471 12903
rect 11241 12903 11299 12909
rect 11241 12900 11253 12903
rect 10413 12863 10471 12869
rect 10796 12872 11253 12900
rect 10796 12841 10824 12872
rect 11241 12869 11253 12872
rect 11287 12900 11299 12903
rect 12066 12900 12072 12912
rect 11287 12872 12072 12900
rect 11287 12869 11299 12872
rect 11241 12863 11299 12869
rect 12066 12860 12072 12872
rect 12124 12860 12130 12912
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 1504 12804 2360 12832
rect 3068 12804 3249 12832
rect 1854 12656 1860 12708
rect 1912 12656 1918 12708
rect 2332 12705 2360 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3421 12835 3479 12841
rect 3421 12801 3433 12835
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 11057 12835 11115 12841
rect 11057 12801 11069 12835
rect 11103 12832 11115 12835
rect 11330 12832 11336 12844
rect 11103 12804 11336 12832
rect 11103 12801 11115 12804
rect 11057 12795 11115 12801
rect 2590 12764 2596 12776
rect 2424 12736 2596 12764
rect 2317 12699 2375 12705
rect 2317 12665 2329 12699
rect 2363 12665 2375 12699
rect 2317 12659 2375 12665
rect 1949 12631 2007 12637
rect 1949 12597 1961 12631
rect 1995 12628 2007 12631
rect 2424 12628 2452 12736
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 2866 12724 2872 12776
rect 2924 12764 2930 12776
rect 3436 12764 3464 12795
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 2924 12736 3464 12764
rect 7101 12767 7159 12773
rect 2924 12724 2930 12736
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 7466 12764 7472 12776
rect 7147 12736 7472 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 9217 12767 9275 12773
rect 9217 12764 9229 12767
rect 7668 12736 9229 12764
rect 7668 12705 7696 12736
rect 9217 12733 9229 12736
rect 9263 12733 9275 12767
rect 9217 12727 9275 12733
rect 9490 12724 9496 12776
rect 9548 12724 9554 12776
rect 11606 12764 11612 12776
rect 10428 12736 11612 12764
rect 7653 12699 7711 12705
rect 7653 12665 7665 12699
rect 7699 12665 7711 12699
rect 7653 12659 7711 12665
rect 1995 12600 2452 12628
rect 2501 12631 2559 12637
rect 1995 12597 2007 12600
rect 1949 12591 2007 12597
rect 2501 12597 2513 12631
rect 2547 12628 2559 12631
rect 2682 12628 2688 12640
rect 2547 12600 2688 12628
rect 2547 12597 2559 12600
rect 2501 12591 2559 12597
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 3234 12588 3240 12640
rect 3292 12588 3298 12640
rect 7466 12588 7472 12640
rect 7524 12588 7530 12640
rect 7742 12588 7748 12640
rect 7800 12588 7806 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10428 12637 10456 12736
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 11716 12764 11744 12795
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 12176 12832 12204 12940
rect 13832 12940 15056 12968
rect 13832 12912 13860 12940
rect 12529 12903 12587 12909
rect 12529 12869 12541 12903
rect 12575 12900 12587 12903
rect 13814 12900 13820 12912
rect 12575 12872 13820 12900
rect 12575 12869 12587 12872
rect 12529 12863 12587 12869
rect 13004 12841 13032 12872
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 14182 12860 14188 12912
rect 14240 12860 14246 12912
rect 14642 12900 14648 12912
rect 14476 12872 14648 12900
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 12176 12804 12357 12832
rect 12345 12801 12357 12804
rect 12391 12832 12403 12835
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12391 12804 12817 12832
rect 12391 12801 12403 12804
rect 12345 12795 12403 12801
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 12989 12835 13047 12841
rect 12989 12801 13001 12835
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13262 12792 13268 12844
rect 13320 12832 13326 12844
rect 14476 12841 14504 12872
rect 14642 12860 14648 12872
rect 14700 12900 14706 12912
rect 14918 12900 14924 12912
rect 14700 12872 14924 12900
rect 14700 12860 14706 12872
rect 14918 12860 14924 12872
rect 14976 12860 14982 12912
rect 13725 12835 13783 12841
rect 13725 12832 13737 12835
rect 13320 12804 13737 12832
rect 13320 12792 13326 12804
rect 13725 12801 13737 12804
rect 13771 12801 13783 12835
rect 13725 12795 13783 12801
rect 13909 12835 13967 12841
rect 13909 12801 13921 12835
rect 13955 12832 13967 12835
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 13955 12804 14381 12832
rect 13955 12801 13967 12804
rect 13909 12795 13967 12801
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 12250 12764 12256 12776
rect 11716 12736 12256 12764
rect 12250 12724 12256 12736
rect 12308 12764 12314 12776
rect 13817 12767 13875 12773
rect 13817 12764 13829 12767
rect 12308 12736 13829 12764
rect 12308 12724 12314 12736
rect 13817 12733 13829 12736
rect 13863 12733 13875 12767
rect 14384 12764 14412 12795
rect 14734 12792 14740 12844
rect 14792 12792 14798 12844
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12832 14887 12835
rect 15028 12832 15056 12940
rect 14875 12804 15056 12832
rect 14875 12801 14887 12804
rect 14829 12795 14887 12801
rect 14921 12767 14979 12773
rect 14921 12764 14933 12767
rect 14384 12736 14933 12764
rect 13817 12727 13875 12733
rect 14921 12733 14933 12736
rect 14967 12733 14979 12767
rect 14921 12727 14979 12733
rect 11330 12656 11336 12708
rect 11388 12696 11394 12708
rect 12069 12699 12127 12705
rect 12069 12696 12081 12699
rect 11388 12668 12081 12696
rect 11388 12656 11394 12668
rect 12069 12665 12081 12668
rect 12115 12665 12127 12699
rect 12069 12659 12127 12665
rect 13262 12656 13268 12708
rect 13320 12696 13326 12708
rect 14645 12699 14703 12705
rect 14645 12696 14657 12699
rect 13320 12668 14657 12696
rect 13320 12656 13326 12668
rect 14645 12665 14657 12668
rect 14691 12665 14703 12699
rect 14645 12659 14703 12665
rect 10229 12631 10287 12637
rect 10229 12628 10241 12631
rect 9824 12600 10241 12628
rect 9824 12588 9830 12600
rect 10229 12597 10241 12600
rect 10275 12597 10287 12631
rect 10229 12591 10287 12597
rect 10413 12631 10471 12637
rect 10413 12597 10425 12631
rect 10459 12597 10471 12631
rect 10413 12591 10471 12597
rect 12710 12588 12716 12640
rect 12768 12588 12774 12640
rect 12894 12588 12900 12640
rect 12952 12588 12958 12640
rect 1104 12538 15456 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 15456 12538
rect 1104 12464 15456 12486
rect 2590 12384 2596 12436
rect 2648 12384 2654 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4706 12424 4712 12436
rect 4295 12396 4712 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 7466 12384 7472 12436
rect 7524 12424 7530 12436
rect 7653 12427 7711 12433
rect 7653 12424 7665 12427
rect 7524 12396 7665 12424
rect 7524 12384 7530 12396
rect 7653 12393 7665 12396
rect 7699 12393 7711 12427
rect 7653 12387 7711 12393
rect 8202 12384 8208 12436
rect 8260 12424 8266 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8260 12396 9045 12424
rect 8260 12384 8266 12396
rect 9033 12393 9045 12396
rect 9079 12393 9091 12427
rect 9033 12387 9091 12393
rect 11606 12384 11612 12436
rect 11664 12384 11670 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 13909 12427 13967 12433
rect 13909 12424 13921 12427
rect 13872 12396 13921 12424
rect 13872 12384 13878 12396
rect 13909 12393 13921 12396
rect 13955 12393 13967 12427
rect 13909 12387 13967 12393
rect 1581 12359 1639 12365
rect 1581 12325 1593 12359
rect 1627 12356 1639 12359
rect 1762 12356 1768 12368
rect 1627 12328 1768 12356
rect 1627 12325 1639 12328
rect 1581 12319 1639 12325
rect 1762 12316 1768 12328
rect 1820 12356 1826 12368
rect 1949 12359 2007 12365
rect 1949 12356 1961 12359
rect 1820 12328 1961 12356
rect 1820 12316 1826 12328
rect 1949 12325 1961 12328
rect 1995 12325 2007 12359
rect 1949 12319 2007 12325
rect 2133 12359 2191 12365
rect 2133 12325 2145 12359
rect 2179 12356 2191 12359
rect 2314 12356 2320 12368
rect 2179 12328 2320 12356
rect 2179 12325 2191 12328
rect 2133 12319 2191 12325
rect 2314 12316 2320 12328
rect 2372 12356 2378 12368
rect 2455 12359 2513 12365
rect 2455 12356 2467 12359
rect 2372 12328 2467 12356
rect 2372 12316 2378 12328
rect 2455 12325 2467 12328
rect 2501 12325 2513 12359
rect 2455 12319 2513 12325
rect 2682 12248 2688 12300
rect 2740 12248 2746 12300
rect 3878 12248 3884 12300
rect 3936 12248 3942 12300
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 5077 12291 5135 12297
rect 5077 12288 5089 12291
rect 4672 12260 5089 12288
rect 4672 12248 4678 12260
rect 5077 12257 5089 12260
rect 5123 12288 5135 12291
rect 5258 12288 5264 12300
rect 5123 12260 5264 12288
rect 5123 12257 5135 12260
rect 5077 12251 5135 12257
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 8754 12288 8760 12300
rect 7116 12260 8760 12288
rect 842 12180 848 12232
rect 900 12220 906 12232
rect 1397 12223 1455 12229
rect 1397 12220 1409 12223
rect 900 12192 1409 12220
rect 900 12180 906 12192
rect 1397 12189 1409 12192
rect 1443 12189 1455 12223
rect 1397 12183 1455 12189
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 3329 12223 3387 12229
rect 3329 12220 3341 12223
rect 2464 12192 3341 12220
rect 2464 12180 2470 12192
rect 3329 12189 3341 12192
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 4525 12223 4583 12229
rect 4525 12220 4537 12223
rect 3476 12192 4537 12220
rect 3476 12180 3482 12192
rect 4525 12189 4537 12192
rect 4571 12220 4583 12223
rect 4709 12223 4767 12229
rect 4571 12192 4660 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 1670 12112 1676 12164
rect 1728 12152 1734 12164
rect 2038 12152 2044 12164
rect 1728 12124 2044 12152
rect 1728 12112 1734 12124
rect 2038 12112 2044 12124
rect 2096 12112 2102 12164
rect 2317 12155 2375 12161
rect 2317 12121 2329 12155
rect 2363 12152 2375 12155
rect 2866 12152 2872 12164
rect 2363 12124 2872 12152
rect 2363 12121 2375 12124
rect 2317 12115 2375 12121
rect 2866 12112 2872 12124
rect 2924 12112 2930 12164
rect 3050 12112 3056 12164
rect 3108 12112 3114 12164
rect 4249 12155 4307 12161
rect 4249 12121 4261 12155
rect 4295 12152 4307 12155
rect 4632 12152 4660 12192
rect 4709 12189 4721 12223
rect 4755 12220 4767 12223
rect 4798 12220 4804 12232
rect 4755 12192 4804 12220
rect 4755 12189 4767 12192
rect 4709 12183 4767 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 4985 12223 5043 12229
rect 4985 12189 4997 12223
rect 5031 12220 5043 12223
rect 6178 12220 6184 12232
rect 5031 12192 6184 12220
rect 5031 12189 5043 12192
rect 4985 12183 5043 12189
rect 6178 12180 6184 12192
rect 6236 12180 6242 12232
rect 6914 12180 6920 12232
rect 6972 12180 6978 12232
rect 7116 12229 7144 12260
rect 8754 12248 8760 12260
rect 8812 12288 8818 12300
rect 9214 12288 9220 12300
rect 8812 12260 9220 12288
rect 8812 12248 8818 12260
rect 9214 12248 9220 12260
rect 9272 12248 9278 12300
rect 13924 12288 13952 12387
rect 14550 12384 14556 12436
rect 14608 12424 14614 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 14608 12396 14933 12424
rect 14608 12384 14614 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 14921 12387 14979 12393
rect 13924 12260 14780 12288
rect 7101 12223 7159 12229
rect 7101 12189 7113 12223
rect 7147 12189 7159 12223
rect 7101 12183 7159 12189
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12220 7435 12223
rect 7466 12220 7472 12232
rect 7423 12192 7472 12220
rect 7423 12189 7435 12192
rect 7377 12183 7435 12189
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 7742 12180 7748 12232
rect 7800 12220 7806 12232
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7800 12192 7849 12220
rect 7800 12180 7806 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 9125 12223 9183 12229
rect 9125 12189 9137 12223
rect 9171 12220 9183 12223
rect 9398 12220 9404 12232
rect 9171 12192 9404 12220
rect 9171 12189 9183 12192
rect 9125 12183 9183 12189
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 9548 12192 11345 12220
rect 9548 12180 9554 12192
rect 11333 12189 11345 12192
rect 11379 12220 11391 12223
rect 12158 12220 12164 12232
rect 11379 12192 12164 12220
rect 11379 12189 11391 12192
rect 11333 12183 11391 12189
rect 12158 12180 12164 12192
rect 12216 12180 12222 12232
rect 14182 12180 14188 12232
rect 14240 12180 14246 12232
rect 14366 12180 14372 12232
rect 14424 12180 14430 12232
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 4893 12155 4951 12161
rect 4893 12152 4905 12155
rect 4295 12124 4568 12152
rect 4632 12124 4905 12152
rect 4295 12121 4307 12124
rect 4249 12115 4307 12121
rect 2774 12044 2780 12096
rect 2832 12084 2838 12096
rect 3145 12087 3203 12093
rect 3145 12084 3157 12087
rect 2832 12056 3157 12084
rect 2832 12044 2838 12056
rect 3145 12053 3157 12056
rect 3191 12053 3203 12087
rect 3145 12047 3203 12053
rect 4430 12044 4436 12096
rect 4488 12044 4494 12096
rect 4540 12093 4568 12124
rect 4893 12121 4905 12124
rect 4939 12121 4951 12155
rect 4893 12115 4951 12121
rect 6825 12155 6883 12161
rect 6825 12121 6837 12155
rect 6871 12152 6883 12155
rect 8938 12152 8944 12164
rect 6871 12124 7788 12152
rect 6871 12121 6883 12124
rect 6825 12115 6883 12121
rect 4525 12087 4583 12093
rect 4525 12053 4537 12087
rect 4571 12053 4583 12087
rect 4525 12047 4583 12053
rect 7101 12087 7159 12093
rect 7101 12053 7113 12087
rect 7147 12084 7159 12087
rect 7190 12084 7196 12096
rect 7147 12056 7196 12084
rect 7147 12053 7159 12056
rect 7101 12047 7159 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 7282 12044 7288 12096
rect 7340 12044 7346 12096
rect 7760 12084 7788 12124
rect 8864 12124 8944 12152
rect 8864 12084 8892 12124
rect 8938 12112 8944 12124
rect 8996 12152 9002 12164
rect 9769 12155 9827 12161
rect 9769 12152 9781 12155
rect 8996 12124 9781 12152
rect 8996 12112 9002 12124
rect 9769 12121 9781 12124
rect 9815 12121 9827 12155
rect 9769 12115 9827 12121
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 11793 12155 11851 12161
rect 11793 12152 11805 12155
rect 11296 12124 11805 12152
rect 11296 12112 11302 12124
rect 11793 12121 11805 12124
rect 11839 12152 11851 12155
rect 11882 12152 11888 12164
rect 11839 12124 11888 12152
rect 11839 12121 11851 12124
rect 11793 12115 11851 12121
rect 11882 12112 11888 12124
rect 11940 12112 11946 12164
rect 11974 12112 11980 12164
rect 12032 12112 12038 12164
rect 12434 12112 12440 12164
rect 12492 12112 12498 12164
rect 13814 12152 13820 12164
rect 13662 12124 13820 12152
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 14274 12112 14280 12164
rect 14332 12152 14338 12164
rect 14476 12152 14504 12183
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 14752 12229 14780 12260
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 14332 12124 14504 12152
rect 14332 12112 14338 12124
rect 7760 12056 8892 12084
rect 1104 11994 15456 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 15456 11994
rect 1104 11920 15456 11942
rect 2225 11883 2283 11889
rect 2225 11849 2237 11883
rect 2271 11880 2283 11883
rect 2866 11880 2872 11892
rect 2271 11852 2872 11880
rect 2271 11849 2283 11852
rect 2225 11843 2283 11849
rect 2866 11840 2872 11852
rect 2924 11840 2930 11892
rect 3878 11840 3884 11892
rect 3936 11880 3942 11892
rect 3973 11883 4031 11889
rect 3973 11880 3985 11883
rect 3936 11852 3985 11880
rect 3936 11840 3942 11852
rect 3973 11849 3985 11852
rect 4019 11849 4031 11883
rect 3973 11843 4031 11849
rect 4430 11840 4436 11892
rect 4488 11880 4494 11892
rect 4488 11852 4752 11880
rect 4488 11840 4494 11852
rect 1762 11772 1768 11824
rect 1820 11772 1826 11824
rect 3234 11812 3240 11824
rect 2516 11784 3240 11812
rect 842 11704 848 11756
rect 900 11744 906 11756
rect 1397 11747 1455 11753
rect 1397 11744 1409 11747
rect 900 11716 1409 11744
rect 900 11704 906 11716
rect 1397 11713 1409 11716
rect 1443 11713 1455 11747
rect 1397 11707 1455 11713
rect 2314 11704 2320 11756
rect 2372 11704 2378 11756
rect 2516 11753 2544 11784
rect 3234 11772 3240 11784
rect 3292 11772 3298 11824
rect 4141 11815 4199 11821
rect 4141 11781 4153 11815
rect 4187 11812 4199 11815
rect 4187 11784 4292 11812
rect 4187 11781 4199 11784
rect 4141 11775 4199 11781
rect 2501 11747 2559 11753
rect 2501 11713 2513 11747
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 2774 11704 2780 11756
rect 2832 11704 2838 11756
rect 3050 11704 3056 11756
rect 3108 11704 3114 11756
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 3234 11676 3240 11688
rect 2639 11648 3240 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 3234 11636 3240 11648
rect 3292 11636 3298 11688
rect 4264 11676 4292 11784
rect 4338 11772 4344 11824
rect 4396 11772 4402 11824
rect 4614 11812 4620 11824
rect 4448 11784 4620 11812
rect 4448 11753 4476 11784
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 4724 11821 4752 11852
rect 6178 11840 6184 11892
rect 6236 11840 6242 11892
rect 7190 11840 7196 11892
rect 7248 11840 7254 11892
rect 9214 11840 9220 11892
rect 9272 11840 9278 11892
rect 11238 11840 11244 11892
rect 11296 11840 11302 11892
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12066 11840 12072 11892
rect 12124 11840 12130 11892
rect 12250 11889 12256 11892
rect 12237 11883 12256 11889
rect 12237 11880 12249 11883
rect 12176 11852 12249 11880
rect 4709 11815 4767 11821
rect 4709 11781 4721 11815
rect 4755 11781 4767 11815
rect 7282 11812 7288 11824
rect 5934 11784 7288 11812
rect 4709 11775 4767 11781
rect 7282 11772 7288 11784
rect 7340 11772 7346 11824
rect 9766 11772 9772 11824
rect 9824 11772 9830 11824
rect 10502 11772 10508 11824
rect 10560 11772 10566 11824
rect 4433 11747 4491 11753
rect 4433 11713 4445 11747
rect 4479 11713 4491 11747
rect 4433 11707 4491 11713
rect 6546 11704 6552 11756
rect 6604 11704 6610 11756
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11744 6883 11747
rect 8662 11744 8668 11756
rect 6871 11716 8668 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 4706 11676 4712 11688
rect 4264 11648 4712 11676
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 2038 11568 2044 11620
rect 2096 11568 2102 11620
rect 2685 11611 2743 11617
rect 2685 11577 2697 11611
rect 2731 11608 2743 11611
rect 3513 11611 3571 11617
rect 3513 11608 3525 11611
rect 2731 11580 3525 11608
rect 2731 11577 2743 11580
rect 2685 11571 2743 11577
rect 3513 11577 3525 11580
rect 3559 11577 3571 11611
rect 3513 11571 3571 11577
rect 5810 11568 5816 11620
rect 5868 11608 5874 11620
rect 6840 11608 6868 11707
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 8754 11704 8760 11756
rect 8812 11744 8818 11756
rect 9125 11747 9183 11753
rect 9125 11744 9137 11747
rect 8812 11716 9137 11744
rect 8812 11704 8818 11716
rect 9125 11713 9137 11716
rect 9171 11713 9183 11747
rect 9125 11707 9183 11713
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11744 11851 11747
rect 12176 11744 12204 11852
rect 12237 11849 12249 11852
rect 12237 11843 12256 11849
rect 12250 11840 12256 11843
rect 12308 11840 12314 11892
rect 12739 11883 12797 11889
rect 12739 11849 12751 11883
rect 12785 11880 12797 11883
rect 12986 11880 12992 11892
rect 12785 11852 12992 11880
rect 12785 11849 12797 11852
rect 12739 11843 12797 11849
rect 12986 11840 12992 11852
rect 13044 11840 13050 11892
rect 13814 11840 13820 11892
rect 13872 11840 13878 11892
rect 14550 11840 14556 11892
rect 14608 11840 14614 11892
rect 12411 11815 12469 11821
rect 12411 11781 12423 11815
rect 12457 11812 12469 11815
rect 12457 11781 12480 11812
rect 12411 11775 12480 11781
rect 12452 11744 12480 11775
rect 12526 11772 12532 11824
rect 12584 11772 12590 11824
rect 11839 11716 12204 11744
rect 12406 11716 12480 11744
rect 13909 11747 13967 11753
rect 11839 11713 11851 11716
rect 11793 11707 11851 11713
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 9490 11676 9496 11688
rect 9088 11648 9496 11676
rect 9088 11636 9094 11648
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 12406 11676 12434 11716
rect 13909 11713 13921 11747
rect 13955 11744 13967 11747
rect 13998 11744 14004 11756
rect 13955 11716 14004 11744
rect 13955 11713 13967 11716
rect 13909 11707 13967 11713
rect 13998 11704 14004 11716
rect 14056 11704 14062 11756
rect 14642 11704 14648 11756
rect 14700 11704 14706 11756
rect 14918 11704 14924 11756
rect 14976 11704 14982 11756
rect 11940 11648 12434 11676
rect 11940 11636 11946 11648
rect 5868 11580 6868 11608
rect 5868 11568 5874 11580
rect 12434 11568 12440 11620
rect 12492 11608 12498 11620
rect 12897 11611 12955 11617
rect 12897 11608 12909 11611
rect 12492 11580 12909 11608
rect 12492 11568 12498 11580
rect 12897 11577 12909 11580
rect 12943 11577 12955 11611
rect 12897 11571 12955 11577
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 2314 11540 2320 11552
rect 1627 11512 2320 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 2314 11500 2320 11512
rect 2372 11500 2378 11552
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 2961 11543 3019 11549
rect 2961 11540 2973 11543
rect 2832 11512 2973 11540
rect 2832 11500 2838 11512
rect 2961 11509 2973 11512
rect 3007 11509 3019 11543
rect 2961 11503 3019 11509
rect 4157 11543 4215 11549
rect 4157 11509 4169 11543
rect 4203 11540 4215 11543
rect 6178 11540 6184 11552
rect 4203 11512 6184 11540
rect 4203 11509 4215 11512
rect 4157 11503 4215 11509
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 6454 11500 6460 11552
rect 6512 11500 6518 11552
rect 7190 11500 7196 11552
rect 7248 11500 7254 11552
rect 7282 11500 7288 11552
rect 7340 11540 7346 11552
rect 7377 11543 7435 11549
rect 7377 11540 7389 11543
rect 7340 11512 7389 11540
rect 7340 11500 7346 11512
rect 7377 11509 7389 11512
rect 7423 11509 7435 11543
rect 7377 11503 7435 11509
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 12253 11543 12311 11549
rect 12253 11540 12265 11543
rect 11756 11512 12265 11540
rect 11756 11500 11762 11512
rect 12253 11509 12265 11512
rect 12299 11509 12311 11543
rect 12253 11503 12311 11509
rect 12710 11500 12716 11552
rect 12768 11500 12774 11552
rect 14366 11500 14372 11552
rect 14424 11540 14430 11552
rect 14829 11543 14887 11549
rect 14829 11540 14841 11543
rect 14424 11512 14841 11540
rect 14424 11500 14430 11512
rect 14829 11509 14841 11512
rect 14875 11509 14887 11543
rect 14829 11503 14887 11509
rect 1104 11450 15456 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 15456 11450
rect 1104 11376 15456 11398
rect 2314 11296 2320 11348
rect 2372 11336 2378 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 2372 11308 3249 11336
rect 2372 11296 2378 11308
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 4246 11336 4252 11348
rect 3237 11299 3295 11305
rect 4080 11308 4252 11336
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11237 1639 11271
rect 3050 11268 3056 11280
rect 1581 11231 1639 11237
rect 2700 11240 3056 11268
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 1596 11132 1624 11231
rect 2700 11209 2728 11240
rect 3050 11228 3056 11240
rect 3108 11228 3114 11280
rect 2685 11203 2743 11209
rect 2685 11169 2697 11203
rect 2731 11169 2743 11203
rect 2685 11163 2743 11169
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3234 11200 3240 11212
rect 2823 11172 3240 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 1596 11104 2973 11132
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3053 11135 3111 11141
rect 3053 11101 3065 11135
rect 3099 11101 3111 11135
rect 3053 11095 3111 11101
rect 3329 11135 3387 11141
rect 3329 11101 3341 11135
rect 3375 11132 3387 11135
rect 3418 11132 3424 11144
rect 3375 11104 3424 11132
rect 3375 11101 3387 11104
rect 3329 11095 3387 11101
rect 2225 10999 2283 11005
rect 2225 10965 2237 10999
rect 2271 10996 2283 10999
rect 2498 10996 2504 11008
rect 2271 10968 2504 10996
rect 2271 10965 2283 10968
rect 2225 10959 2283 10965
rect 2498 10956 2504 10968
rect 2556 10956 2562 11008
rect 2976 10996 3004 11095
rect 3068 11064 3096 11095
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 4080 11141 4108 11308
rect 4246 11296 4252 11308
rect 4304 11336 4310 11348
rect 4890 11336 4896 11348
rect 4304 11308 4896 11336
rect 4304 11296 4310 11308
rect 4890 11296 4896 11308
rect 4948 11336 4954 11348
rect 6825 11339 6883 11345
rect 6825 11336 6837 11339
rect 4948 11308 6837 11336
rect 4948 11296 4954 11308
rect 6825 11305 6837 11308
rect 6871 11305 6883 11339
rect 6825 11299 6883 11305
rect 8754 11296 8760 11348
rect 8812 11296 8818 11348
rect 10502 11296 10508 11348
rect 10560 11296 10566 11348
rect 13541 11339 13599 11345
rect 13541 11305 13553 11339
rect 13587 11336 13599 11339
rect 13998 11336 14004 11348
rect 13587 11308 14004 11336
rect 13587 11305 13599 11308
rect 13541 11299 13599 11305
rect 4614 11228 4620 11280
rect 4672 11268 4678 11280
rect 4672 11240 5120 11268
rect 4672 11228 4678 11240
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 4798 11200 4804 11212
rect 4203 11172 4804 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 3605 11135 3663 11141
rect 3605 11101 3617 11135
rect 3651 11132 3663 11135
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3651 11104 4077 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 4249 11135 4307 11141
rect 4249 11101 4261 11135
rect 4295 11101 4307 11135
rect 4249 11095 4307 11101
rect 3513 11067 3571 11073
rect 3513 11064 3525 11067
rect 3068 11036 3525 11064
rect 3513 11033 3525 11036
rect 3559 11033 3571 11067
rect 4264 11064 4292 11095
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 4540 11141 4568 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 5092 11209 5120 11240
rect 5077 11203 5135 11209
rect 5077 11169 5089 11203
rect 5123 11200 5135 11203
rect 5123 11172 7052 11200
rect 5123 11169 5135 11172
rect 5077 11163 5135 11169
rect 7024 11144 7052 11172
rect 7282 11160 7288 11212
rect 7340 11160 7346 11212
rect 13556 11200 13584 11299
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 14918 11296 14924 11348
rect 14976 11296 14982 11348
rect 10428 11172 13584 11200
rect 10428 11144 10456 11172
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 4890 11132 4896 11144
rect 4755 11104 4896 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 4632 11064 4660 11095
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 6454 11092 6460 11144
rect 6512 11092 6518 11144
rect 7006 11092 7012 11144
rect 7064 11092 7070 11144
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11132 9183 11135
rect 9306 11132 9312 11144
rect 9171 11104 9312 11132
rect 9171 11101 9183 11104
rect 9125 11095 9183 11101
rect 9306 11092 9312 11104
rect 9364 11092 9370 11144
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 10410 11132 10416 11144
rect 9456 11104 10416 11132
rect 9456 11092 9462 11104
rect 10410 11092 10416 11104
rect 10468 11092 10474 11144
rect 11790 11092 11796 11144
rect 11848 11132 11854 11144
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 11848 11104 11897 11132
rect 11848 11092 11854 11104
rect 11885 11101 11897 11104
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 11974 11092 11980 11144
rect 12032 11092 12038 11144
rect 12066 11092 12072 11144
rect 12124 11092 12130 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12250 11132 12256 11144
rect 12207 11104 12256 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 14016 11132 14044 11296
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 14016 11104 14289 11132
rect 14277 11101 14289 11104
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14829 11135 14887 11141
rect 14829 11101 14841 11135
rect 14875 11101 14887 11135
rect 14829 11095 14887 11101
rect 4798 11064 4804 11076
rect 4264 11036 4804 11064
rect 3513 11027 3571 11033
rect 4798 11024 4804 11036
rect 4856 11024 4862 11076
rect 4985 11067 5043 11073
rect 4985 11033 4997 11067
rect 5031 11064 5043 11067
rect 5353 11067 5411 11073
rect 5353 11064 5365 11067
rect 5031 11036 5365 11064
rect 5031 11033 5043 11036
rect 4985 11027 5043 11033
rect 5353 11033 5365 11036
rect 5399 11033 5411 11067
rect 9033 11067 9091 11073
rect 9033 11064 9045 11067
rect 8510 11036 9045 11064
rect 5353 11027 5411 11033
rect 9033 11033 9045 11036
rect 9079 11033 9091 11067
rect 9033 11027 9091 11033
rect 13630 11024 13636 11076
rect 13688 11024 13694 11076
rect 14182 11024 14188 11076
rect 14240 11024 14246 11076
rect 14844 11064 14872 11095
rect 15102 11092 15108 11144
rect 15160 11092 15166 11144
rect 15194 11064 15200 11076
rect 14844 11036 15200 11064
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 3878 10996 3884 11008
rect 2976 10968 3884 10996
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 11701 10999 11759 11005
rect 11701 10965 11713 10999
rect 11747 10996 11759 10999
rect 11882 10996 11888 11008
rect 11747 10968 11888 10996
rect 11747 10965 11759 10968
rect 11701 10959 11759 10965
rect 11882 10956 11888 10968
rect 11940 10956 11946 11008
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 14274 10996 14280 11008
rect 12308 10968 14280 10996
rect 12308 10956 12314 10968
rect 14274 10956 14280 10968
rect 14332 10956 14338 11008
rect 14645 10999 14703 11005
rect 14645 10965 14657 10999
rect 14691 10996 14703 10999
rect 14734 10996 14740 11008
rect 14691 10968 14740 10996
rect 14691 10965 14703 10968
rect 14645 10959 14703 10965
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 1104 10906 15456 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 15456 10906
rect 1104 10832 15456 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 2593 10795 2651 10801
rect 2593 10761 2605 10795
rect 2639 10792 2651 10795
rect 4706 10792 4712 10804
rect 2639 10764 4712 10792
rect 2639 10761 2651 10764
rect 2593 10755 2651 10761
rect 1596 10724 1624 10755
rect 4706 10752 4712 10764
rect 4764 10752 4770 10804
rect 6454 10752 6460 10804
rect 6512 10752 6518 10804
rect 9937 10795 9995 10801
rect 9937 10761 9949 10795
rect 9983 10792 9995 10795
rect 10505 10795 10563 10801
rect 10505 10792 10517 10795
rect 9983 10764 10517 10792
rect 9983 10761 9995 10764
rect 9937 10755 9995 10761
rect 10505 10761 10517 10764
rect 10551 10761 10563 10795
rect 12526 10792 12532 10804
rect 10505 10755 10563 10761
rect 12406 10764 12532 10792
rect 4062 10724 4068 10736
rect 1596 10696 4068 10724
rect 4062 10684 4068 10696
rect 4120 10684 4126 10736
rect 4246 10684 4252 10736
rect 4304 10684 4310 10736
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 11885 10727 11943 10733
rect 11885 10724 11897 10727
rect 10192 10696 11897 10724
rect 10192 10684 10198 10696
rect 11885 10693 11897 10696
rect 11931 10724 11943 10727
rect 12406 10724 12434 10764
rect 12526 10752 12532 10764
rect 12584 10752 12590 10804
rect 14182 10724 14188 10736
rect 11931 10696 12434 10724
rect 13662 10696 14188 10724
rect 11931 10693 11943 10696
rect 11885 10687 11943 10693
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 14366 10684 14372 10736
rect 14424 10684 14430 10736
rect 14458 10684 14464 10736
rect 14516 10724 14522 10736
rect 14829 10727 14887 10733
rect 14829 10724 14841 10727
rect 14516 10696 14841 10724
rect 14516 10684 14522 10696
rect 14829 10693 14841 10696
rect 14875 10693 14887 10727
rect 14829 10687 14887 10693
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 900 10628 1409 10656
rect 900 10616 906 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 2498 10616 2504 10668
rect 2556 10616 2562 10668
rect 2685 10659 2743 10665
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 2866 10656 2872 10668
rect 2731 10628 2872 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 2866 10616 2872 10628
rect 2924 10656 2930 10668
rect 5261 10659 5319 10665
rect 2924 10628 3372 10656
rect 2924 10616 2930 10628
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 3234 10588 3240 10600
rect 2823 10560 3240 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 3344 10597 3372 10628
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5994 10656 6000 10668
rect 5307 10628 6000 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5994 10616 6000 10628
rect 6052 10656 6058 10668
rect 6549 10659 6607 10665
rect 6549 10656 6561 10659
rect 6052 10628 6561 10656
rect 6052 10616 6058 10628
rect 6549 10625 6561 10628
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7282 10656 7288 10668
rect 7147 10628 7288 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 3329 10591 3387 10597
rect 3329 10557 3341 10591
rect 3375 10557 3387 10591
rect 6564 10588 6592 10619
rect 7282 10616 7288 10628
rect 7340 10616 7346 10668
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 10502 10616 10508 10668
rect 10560 10616 10566 10668
rect 10689 10659 10747 10665
rect 10689 10625 10701 10659
rect 10735 10656 10747 10659
rect 11238 10656 11244 10668
rect 10735 10628 11244 10656
rect 10735 10625 10747 10628
rect 10689 10619 10747 10625
rect 11238 10616 11244 10628
rect 11296 10616 11302 10668
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10656 11575 10659
rect 11698 10656 11704 10668
rect 11563 10628 11704 10656
rect 11563 10625 11575 10628
rect 11517 10619 11575 10625
rect 11698 10616 11704 10628
rect 11756 10616 11762 10668
rect 12158 10616 12164 10668
rect 12216 10616 12222 10668
rect 14274 10656 14280 10668
rect 13924 10628 14280 10656
rect 7466 10588 7472 10600
rect 6564 10560 7472 10588
rect 3329 10551 3387 10557
rect 7466 10548 7472 10560
rect 7524 10588 7530 10600
rect 9398 10588 9404 10600
rect 7524 10560 9404 10588
rect 7524 10548 7530 10560
rect 9398 10548 9404 10560
rect 9456 10548 9462 10600
rect 13924 10597 13952 10628
rect 14274 10616 14280 10628
rect 14332 10616 14338 10668
rect 14642 10616 14648 10668
rect 14700 10616 14706 10668
rect 14734 10616 14740 10668
rect 14792 10616 14798 10668
rect 12437 10591 12495 10597
rect 12437 10588 12449 10591
rect 12084 10560 12449 10588
rect 3050 10480 3056 10532
rect 3108 10520 3114 10532
rect 3421 10523 3479 10529
rect 3421 10520 3433 10523
rect 3108 10492 3433 10520
rect 3108 10480 3114 10492
rect 3421 10489 3433 10492
rect 3467 10489 3479 10523
rect 3421 10483 3479 10489
rect 3878 10480 3884 10532
rect 3936 10480 3942 10532
rect 12084 10529 12112 10560
rect 12437 10557 12449 10560
rect 12483 10557 12495 10591
rect 12437 10551 12495 10557
rect 13909 10591 13967 10597
rect 13909 10557 13921 10591
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 12069 10523 12127 10529
rect 12069 10489 12081 10523
rect 12115 10489 12127 10523
rect 12069 10483 12127 10489
rect 3142 10412 3148 10464
rect 3200 10412 3206 10464
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 3786 10452 3792 10464
rect 3283 10424 3792 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 3786 10412 3792 10424
rect 3844 10412 3850 10464
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 5353 10455 5411 10461
rect 5353 10452 5365 10455
rect 5316 10424 5365 10452
rect 5316 10412 5322 10424
rect 5353 10421 5365 10424
rect 5399 10421 5411 10455
rect 5353 10415 5411 10421
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7009 10455 7067 10461
rect 7009 10452 7021 10455
rect 6972 10424 7021 10452
rect 6972 10412 6978 10424
rect 7009 10421 7021 10424
rect 7055 10421 7067 10455
rect 7009 10415 7067 10421
rect 9306 10412 9312 10464
rect 9364 10452 9370 10464
rect 9769 10455 9827 10461
rect 9769 10452 9781 10455
rect 9364 10424 9781 10452
rect 9364 10412 9370 10424
rect 9769 10421 9781 10424
rect 9815 10421 9827 10455
rect 9769 10415 9827 10421
rect 9950 10412 9956 10464
rect 10008 10412 10014 10464
rect 10318 10412 10324 10464
rect 10376 10412 10382 10464
rect 11882 10412 11888 10464
rect 11940 10412 11946 10464
rect 13998 10412 14004 10464
rect 14056 10452 14062 10464
rect 14093 10455 14151 10461
rect 14093 10452 14105 10455
rect 14056 10424 14105 10452
rect 14056 10412 14062 10424
rect 14093 10421 14105 10424
rect 14139 10421 14151 10455
rect 14093 10415 14151 10421
rect 1104 10362 15456 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 15456 10362
rect 1104 10288 15456 10310
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10873 10251 10931 10257
rect 10873 10248 10885 10251
rect 10008 10220 10885 10248
rect 10008 10208 10014 10220
rect 10873 10217 10885 10220
rect 10919 10217 10931 10251
rect 10873 10211 10931 10217
rect 11698 10208 11704 10260
rect 11756 10208 11762 10260
rect 12066 10208 12072 10260
rect 12124 10248 12130 10260
rect 12124 10220 12388 10248
rect 12124 10208 12130 10220
rect 1857 10183 1915 10189
rect 1857 10149 1869 10183
rect 1903 10180 1915 10183
rect 2038 10180 2044 10192
rect 1903 10152 2044 10180
rect 1903 10149 1915 10152
rect 1857 10143 1915 10149
rect 2038 10140 2044 10152
rect 2096 10140 2102 10192
rect 5626 10140 5632 10192
rect 5684 10180 5690 10192
rect 5997 10183 6055 10189
rect 5997 10180 6009 10183
rect 5684 10152 6009 10180
rect 5684 10140 5690 10152
rect 5997 10149 6009 10152
rect 6043 10149 6055 10183
rect 5997 10143 6055 10149
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 12032 10152 12204 10180
rect 12032 10140 12038 10152
rect 4249 10115 4307 10121
rect 4249 10081 4261 10115
rect 4295 10112 4307 10115
rect 4614 10112 4620 10124
rect 4295 10084 4620 10112
rect 4295 10081 4307 10084
rect 4249 10075 4307 10081
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 5592 10084 6316 10112
rect 5592 10072 5598 10084
rect 2222 10004 2228 10056
rect 2280 10004 2286 10056
rect 6288 10053 6316 10084
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 8757 10115 8815 10121
rect 8757 10112 8769 10115
rect 7340 10084 8769 10112
rect 7340 10072 7346 10084
rect 8757 10081 8769 10084
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 9030 10072 9036 10124
rect 9088 10072 9094 10124
rect 9306 10072 9312 10124
rect 9364 10072 9370 10124
rect 10502 10072 10508 10124
rect 10560 10112 10566 10124
rect 10781 10115 10839 10121
rect 10781 10112 10793 10115
rect 10560 10084 10793 10112
rect 10560 10072 10566 10084
rect 10781 10081 10793 10084
rect 10827 10112 10839 10115
rect 12066 10112 12072 10124
rect 10827 10084 12072 10112
rect 10827 10081 10839 10084
rect 10781 10075 10839 10081
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 6362 10044 6368 10056
rect 6319 10016 6368 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 1489 9979 1547 9985
rect 1489 9945 1501 9979
rect 1535 9976 1547 9979
rect 1762 9976 1768 9988
rect 1535 9948 1768 9976
rect 1535 9945 1547 9948
rect 1489 9939 1547 9945
rect 1762 9936 1768 9948
rect 1820 9976 1826 9988
rect 4525 9979 4583 9985
rect 1820 9948 2084 9976
rect 1820 9936 1826 9948
rect 1946 9868 1952 9920
rect 2004 9868 2010 9920
rect 2056 9917 2084 9948
rect 4525 9945 4537 9979
rect 4571 9976 4583 9979
rect 4614 9976 4620 9988
rect 4571 9948 4620 9976
rect 4571 9945 4583 9948
rect 4525 9939 4583 9945
rect 4614 9936 4620 9948
rect 4672 9936 4678 9988
rect 5258 9936 5264 9988
rect 5316 9936 5322 9988
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9877 2099 9911
rect 6472 9908 6500 10007
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 6822 10044 6828 10056
rect 6687 10016 6828 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 7006 10004 7012 10056
rect 7064 10004 7070 10056
rect 11057 10047 11115 10053
rect 11057 10013 11069 10047
rect 11103 10044 11115 10047
rect 11164 10044 11192 10084
rect 12066 10072 12072 10084
rect 12124 10072 12130 10124
rect 12176 10112 12204 10152
rect 12250 10140 12256 10192
rect 12308 10140 12314 10192
rect 12360 10180 12388 10220
rect 13446 10208 13452 10260
rect 13504 10208 13510 10260
rect 14553 10251 14611 10257
rect 14553 10217 14565 10251
rect 14599 10248 14611 10251
rect 14642 10248 14648 10260
rect 14599 10220 14648 10248
rect 14599 10217 14611 10220
rect 14553 10211 14611 10217
rect 14568 10180 14596 10211
rect 14642 10208 14648 10220
rect 14700 10208 14706 10260
rect 12360 10152 14596 10180
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 12176 10084 12725 10112
rect 12713 10081 12725 10084
rect 12759 10081 12771 10115
rect 13998 10112 14004 10124
rect 12713 10075 12771 10081
rect 13648 10084 14004 10112
rect 11103 10016 11192 10044
rect 11103 10013 11115 10016
rect 11057 10007 11115 10013
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 13648 10053 13676 10084
rect 13998 10072 14004 10084
rect 14056 10072 14062 10124
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 11296 10016 12357 10044
rect 11296 10004 11302 10016
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12345 10007 12403 10013
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10013 12587 10047
rect 12529 10007 12587 10013
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 13909 10047 13967 10053
rect 13909 10013 13921 10047
rect 13955 10044 13967 10047
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13955 10016 14105 10044
rect 13955 10013 13967 10016
rect 13909 10007 13967 10013
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 6917 9979 6975 9985
rect 6917 9945 6929 9979
rect 6963 9976 6975 9979
rect 7285 9979 7343 9985
rect 7285 9976 7297 9979
rect 6963 9948 7297 9976
rect 6963 9945 6975 9948
rect 6917 9939 6975 9945
rect 7285 9945 7297 9948
rect 7331 9945 7343 9979
rect 9306 9976 9312 9988
rect 8510 9948 9312 9976
rect 7285 9939 7343 9945
rect 9306 9936 9312 9948
rect 9364 9936 9370 9988
rect 10318 9936 10324 9988
rect 10376 9936 10382 9988
rect 11790 9936 11796 9988
rect 11848 9976 11854 9988
rect 11885 9979 11943 9985
rect 11885 9976 11897 9979
rect 11848 9948 11897 9976
rect 11848 9936 11854 9948
rect 11885 9945 11897 9948
rect 11931 9976 11943 9979
rect 12250 9976 12256 9988
rect 11931 9948 12256 9976
rect 11931 9945 11943 9948
rect 11885 9939 11943 9945
rect 12250 9936 12256 9948
rect 12308 9976 12314 9988
rect 12308 9948 12434 9976
rect 12308 9936 12314 9948
rect 7098 9908 7104 9920
rect 6472 9880 7104 9908
rect 2041 9871 2099 9877
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 11974 9908 11980 9920
rect 11112 9880 11980 9908
rect 11112 9868 11118 9880
rect 11974 9868 11980 9880
rect 12032 9868 12038 9920
rect 12066 9868 12072 9920
rect 12124 9868 12130 9920
rect 12406 9908 12434 9948
rect 12544 9908 12572 10007
rect 14274 10004 14280 10056
rect 14332 10004 14338 10056
rect 14369 10047 14427 10053
rect 14369 10013 14381 10047
rect 14415 10013 14427 10047
rect 14369 10007 14427 10013
rect 14182 9936 14188 9988
rect 14240 9976 14246 9988
rect 14384 9976 14412 10007
rect 14458 10004 14464 10056
rect 14516 10044 14522 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 14516 10016 14657 10044
rect 14516 10004 14522 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 15102 10004 15108 10056
rect 15160 10004 15166 10056
rect 14240 9948 14412 9976
rect 14240 9936 14246 9948
rect 12406 9880 12572 9908
rect 13814 9868 13820 9920
rect 13872 9868 13878 9920
rect 14918 9868 14924 9920
rect 14976 9868 14982 9920
rect 1104 9818 15456 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 15456 9818
rect 1104 9744 15456 9766
rect 2777 9707 2835 9713
rect 2777 9673 2789 9707
rect 2823 9704 2835 9707
rect 2823 9676 3464 9704
rect 2823 9673 2835 9676
rect 2777 9667 2835 9673
rect 2746 9608 3372 9636
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9568 1547 9571
rect 2038 9568 2044 9580
rect 1535 9540 2044 9568
rect 1535 9537 1547 9540
rect 1489 9531 1547 9537
rect 2038 9528 2044 9540
rect 2096 9528 2102 9580
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9537 2283 9571
rect 2225 9531 2283 9537
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2240 9500 2268 9531
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 2746 9568 2774 9608
rect 2556 9540 2774 9568
rect 2556 9528 2562 9540
rect 3050 9528 3056 9580
rect 3108 9528 3114 9580
rect 3344 9577 3372 9608
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9537 3203 9571
rect 3145 9531 3203 9537
rect 3329 9571 3387 9577
rect 3329 9537 3341 9571
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 1995 9472 2268 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 2314 9460 2320 9512
rect 2372 9460 2378 9512
rect 2774 9460 2780 9512
rect 2832 9460 2838 9512
rect 1762 9392 1768 9444
rect 1820 9392 1826 9444
rect 3160 9432 3188 9531
rect 3436 9500 3464 9676
rect 4614 9664 4620 9716
rect 4672 9704 4678 9716
rect 4709 9707 4767 9713
rect 4709 9704 4721 9707
rect 4672 9676 4721 9704
rect 4672 9664 4678 9676
rect 4709 9673 4721 9676
rect 4755 9673 4767 9707
rect 4709 9667 4767 9673
rect 4801 9707 4859 9713
rect 4801 9673 4813 9707
rect 4847 9673 4859 9707
rect 4801 9667 4859 9673
rect 11977 9707 12035 9713
rect 11977 9673 11989 9707
rect 12023 9704 12035 9707
rect 12526 9704 12532 9716
rect 12023 9676 12532 9704
rect 12023 9673 12035 9676
rect 11977 9667 12035 9673
rect 4525 9639 4583 9645
rect 4525 9605 4537 9639
rect 4571 9636 4583 9639
rect 4816 9636 4844 9667
rect 12526 9664 12532 9676
rect 12584 9664 12590 9716
rect 14274 9664 14280 9716
rect 14332 9704 14338 9716
rect 14553 9707 14611 9713
rect 14553 9704 14565 9707
rect 14332 9676 14565 9704
rect 14332 9664 14338 9676
rect 14553 9673 14565 9676
rect 14599 9673 14611 9707
rect 14553 9667 14611 9673
rect 7282 9636 7288 9648
rect 4571 9608 4844 9636
rect 5092 9608 7288 9636
rect 4571 9605 4583 9608
rect 4525 9599 4583 9605
rect 3970 9528 3976 9580
rect 4028 9568 4034 9580
rect 4028 9566 4752 9568
rect 4890 9566 4896 9580
rect 4028 9540 4896 9566
rect 4028 9528 4034 9540
rect 4724 9538 4896 9540
rect 4890 9528 4896 9538
rect 4948 9568 4954 9580
rect 5092 9577 5120 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 7374 9596 7380 9648
rect 7432 9596 7438 9648
rect 8938 9596 8944 9648
rect 8996 9596 9002 9648
rect 9306 9596 9312 9648
rect 9364 9596 9370 9648
rect 10134 9596 10140 9648
rect 10192 9596 10198 9648
rect 14458 9636 14464 9648
rect 12452 9608 14464 9636
rect 5077 9571 5135 9577
rect 5077 9568 5089 9571
rect 4948 9540 5089 9568
rect 4948 9528 4954 9540
rect 5077 9537 5089 9540
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9568 5319 9571
rect 5626 9568 5632 9580
rect 5307 9540 5632 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 6454 9528 6460 9580
rect 6512 9528 6518 9580
rect 9398 9528 9404 9580
rect 9456 9528 9462 9580
rect 10502 9528 10508 9580
rect 10560 9528 10566 9580
rect 10870 9528 10876 9580
rect 10928 9568 10934 9580
rect 10965 9571 11023 9577
rect 10965 9568 10977 9571
rect 10928 9540 10977 9568
rect 10928 9528 10934 9540
rect 10965 9537 10977 9540
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 11149 9571 11207 9577
rect 11149 9537 11161 9571
rect 11195 9537 11207 9571
rect 11149 9531 11207 9537
rect 3436 9472 4936 9500
rect 2240 9404 3188 9432
rect 4157 9435 4215 9441
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 2240 9373 2268 9404
rect 4157 9401 4169 9435
rect 4203 9432 4215 9435
rect 4614 9432 4620 9444
rect 4203 9404 4620 9432
rect 4203 9401 4215 9404
rect 4157 9395 4215 9401
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 4908 9432 4936 9472
rect 4982 9460 4988 9512
rect 5040 9460 5046 9512
rect 5166 9460 5172 9512
rect 5224 9460 5230 9512
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 7190 9500 7196 9512
rect 6779 9472 7196 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 6270 9432 6276 9444
rect 4908 9404 6276 9432
rect 6270 9392 6276 9404
rect 6328 9392 6334 9444
rect 2225 9367 2283 9373
rect 2225 9364 2237 9367
rect 2004 9336 2237 9364
rect 2004 9324 2010 9336
rect 2225 9333 2237 9336
rect 2271 9333 2283 9367
rect 2225 9327 2283 9333
rect 2685 9367 2743 9373
rect 2685 9333 2697 9367
rect 2731 9364 2743 9367
rect 2774 9364 2780 9376
rect 2731 9336 2780 9364
rect 2731 9333 2743 9336
rect 2685 9327 2743 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 3142 9324 3148 9376
rect 3200 9324 3206 9376
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 6748 9364 6776 9463
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 11164 9500 11192 9531
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11296 9540 11621 9568
rect 11296 9528 11302 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 12250 9528 12256 9580
rect 12308 9528 12314 9580
rect 12342 9528 12348 9580
rect 12400 9568 12406 9580
rect 12452 9577 12480 9608
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 12437 9571 12495 9577
rect 12437 9568 12449 9571
rect 12400 9540 12449 9568
rect 12400 9528 12406 9540
rect 12437 9537 12449 9540
rect 12483 9537 12495 9571
rect 12437 9531 12495 9537
rect 13173 9571 13231 9577
rect 13173 9537 13185 9571
rect 13219 9568 13231 9571
rect 13446 9568 13452 9580
rect 13219 9540 13452 9568
rect 13219 9537 13231 9540
rect 13173 9531 13231 9537
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 14642 9528 14648 9580
rect 14700 9528 14706 9580
rect 14918 9528 14924 9580
rect 14976 9528 14982 9580
rect 11422 9500 11428 9512
rect 11164 9472 11428 9500
rect 11422 9460 11428 9472
rect 11480 9460 11486 9512
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 12621 9503 12679 9509
rect 12621 9500 12633 9503
rect 11940 9472 12633 9500
rect 11940 9460 11946 9472
rect 12621 9469 12633 9472
rect 12667 9500 12679 9503
rect 14182 9500 14188 9512
rect 12667 9472 14188 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 14182 9460 14188 9472
rect 14240 9460 14246 9512
rect 12161 9435 12219 9441
rect 12161 9401 12173 9435
rect 12207 9432 12219 9435
rect 12434 9432 12440 9444
rect 12207 9404 12440 9432
rect 12207 9401 12219 9404
rect 12161 9395 12219 9401
rect 12434 9392 12440 9404
rect 12492 9392 12498 9444
rect 4571 9336 6776 9364
rect 11057 9367 11115 9373
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 11057 9333 11069 9367
rect 11103 9364 11115 9367
rect 11514 9364 11520 9376
rect 11103 9336 11520 9364
rect 11103 9333 11115 9336
rect 11057 9327 11115 9333
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 12066 9364 12072 9376
rect 12023 9336 12072 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 13170 9324 13176 9376
rect 13228 9364 13234 9376
rect 13265 9367 13323 9373
rect 13265 9364 13277 9367
rect 13228 9336 13277 9364
rect 13228 9324 13234 9336
rect 13265 9333 13277 9336
rect 13311 9333 13323 9367
rect 13265 9327 13323 9333
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 13412 9336 14841 9364
rect 13412 9324 13418 9336
rect 14829 9333 14841 9336
rect 14875 9333 14887 9367
rect 14829 9327 14887 9333
rect 1104 9274 15456 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 15456 9274
rect 1104 9200 15456 9222
rect 2225 9163 2283 9169
rect 2225 9129 2237 9163
rect 2271 9160 2283 9163
rect 2498 9160 2504 9172
rect 2271 9132 2504 9160
rect 2271 9129 2283 9132
rect 2225 9123 2283 9129
rect 2498 9120 2504 9132
rect 2556 9120 2562 9172
rect 2608 9132 2912 9160
rect 2130 9052 2136 9104
rect 2188 9092 2194 9104
rect 2608 9092 2636 9132
rect 2188 9064 2636 9092
rect 2685 9095 2743 9101
rect 2188 9052 2194 9064
rect 2685 9061 2697 9095
rect 2731 9092 2743 9095
rect 2774 9092 2780 9104
rect 2731 9064 2780 9092
rect 2731 9061 2743 9064
rect 2685 9055 2743 9061
rect 2774 9052 2780 9064
rect 2832 9052 2838 9104
rect 2884 9092 2912 9132
rect 2958 9120 2964 9172
rect 3016 9120 3022 9172
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 4798 9160 4804 9172
rect 4672 9132 4804 9160
rect 4672 9120 4678 9132
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 6420 9132 9076 9160
rect 6420 9120 6426 9132
rect 2884 9064 4384 9092
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 3142 9024 3148 9036
rect 2547 8996 3148 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 3142 8984 3148 8996
rect 3200 8984 3206 9036
rect 842 8916 848 8968
rect 900 8956 906 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 900 8928 1409 8956
rect 900 8916 906 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 2314 8916 2320 8968
rect 2372 8916 2378 8968
rect 2593 8959 2651 8965
rect 2593 8925 2605 8959
rect 2639 8956 2651 8959
rect 2682 8956 2688 8968
rect 2639 8928 2688 8956
rect 2639 8925 2651 8928
rect 2593 8919 2651 8925
rect 2682 8916 2688 8928
rect 2740 8916 2746 8968
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8956 2835 8959
rect 2866 8956 2872 8968
rect 2823 8928 2872 8956
rect 2823 8925 2835 8928
rect 2777 8919 2835 8925
rect 2866 8916 2872 8928
rect 2924 8956 2930 8968
rect 3326 8956 3332 8968
rect 2924 8928 3332 8956
rect 2924 8916 2930 8928
rect 3326 8916 3332 8928
rect 3384 8916 3390 8968
rect 1765 8891 1823 8897
rect 1765 8857 1777 8891
rect 1811 8857 1823 8891
rect 4356 8888 4384 9064
rect 5074 9052 5080 9104
rect 5132 9092 5138 9104
rect 9048 9101 9076 9132
rect 12066 9120 12072 9172
rect 12124 9120 12130 9172
rect 13446 9160 13452 9172
rect 12176 9132 13452 9160
rect 9033 9095 9091 9101
rect 5132 9064 5948 9092
rect 5132 9052 5138 9064
rect 4617 9027 4675 9033
rect 4617 8993 4629 9027
rect 4663 9024 4675 9027
rect 4798 9024 4804 9036
rect 4663 8996 4804 9024
rect 4663 8993 4675 8996
rect 4617 8987 4675 8993
rect 4798 8984 4804 8996
rect 4856 8984 4862 9036
rect 4982 8984 4988 9036
rect 5040 9024 5046 9036
rect 5350 9024 5356 9036
rect 5040 8996 5356 9024
rect 5040 8984 5046 8996
rect 5350 8984 5356 8996
rect 5408 9024 5414 9036
rect 5408 8996 5856 9024
rect 5408 8984 5414 8996
rect 4890 8916 4896 8968
rect 4948 8916 4954 8968
rect 5534 8916 5540 8968
rect 5592 8916 5598 8968
rect 5718 8916 5724 8968
rect 5776 8916 5782 8968
rect 5828 8965 5856 8996
rect 5920 8965 5948 9064
rect 9033 9061 9045 9095
rect 9079 9061 9091 9095
rect 9033 9055 9091 9061
rect 6273 9027 6331 9033
rect 6273 8993 6285 9027
rect 6319 9024 6331 9027
rect 7006 9024 7012 9036
rect 6319 8996 7012 9024
rect 6319 8993 6331 8996
rect 6273 8987 6331 8993
rect 7006 8984 7012 8996
rect 7064 8984 7070 9036
rect 9048 9024 9076 9055
rect 9398 9052 9404 9104
rect 9456 9092 9462 9104
rect 12176 9092 12204 9132
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 14642 9120 14648 9172
rect 14700 9160 14706 9172
rect 14921 9163 14979 9169
rect 14921 9160 14933 9163
rect 14700 9132 14933 9160
rect 14700 9120 14706 9132
rect 14921 9129 14933 9132
rect 14967 9129 14979 9163
rect 14921 9123 14979 9129
rect 9456 9064 12204 9092
rect 9456 9052 9462 9064
rect 10502 9024 10508 9036
rect 9048 8996 10508 9024
rect 10502 8984 10508 8996
rect 10560 9024 10566 9036
rect 10560 8996 10824 9024
rect 10560 8984 10566 8996
rect 5813 8959 5871 8965
rect 5813 8925 5825 8959
rect 5859 8925 5871 8959
rect 5813 8919 5871 8925
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8925 5963 8959
rect 5905 8919 5963 8925
rect 4985 8891 5043 8897
rect 4985 8888 4997 8891
rect 4356 8860 4997 8888
rect 1765 8851 1823 8857
rect 4985 8857 4997 8860
rect 5031 8888 5043 8891
rect 5626 8888 5632 8900
rect 5031 8860 5632 8888
rect 5031 8857 5043 8860
rect 4985 8851 5043 8857
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1780 8820 1808 8851
rect 5626 8848 5632 8860
rect 5684 8848 5690 8900
rect 1854 8820 1860 8832
rect 1627 8792 1860 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1854 8780 1860 8792
rect 1912 8780 1918 8832
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 3970 8820 3976 8832
rect 2096 8792 3976 8820
rect 2096 8780 2102 8792
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4580 8792 4813 8820
rect 4580 8780 4586 8792
rect 4801 8789 4813 8792
rect 4847 8820 4859 8823
rect 5074 8820 5080 8832
rect 4847 8792 5080 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5169 8823 5227 8829
rect 5169 8789 5181 8823
rect 5215 8820 5227 8823
rect 5258 8820 5264 8832
rect 5215 8792 5264 8820
rect 5215 8789 5227 8792
rect 5169 8783 5227 8789
rect 5258 8780 5264 8792
rect 5316 8780 5322 8832
rect 5920 8820 5948 8919
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8536 8928 8953 8956
rect 8536 8916 8542 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 8941 8919 8999 8925
rect 9585 8959 9643 8965
rect 9585 8925 9597 8959
rect 9631 8956 9643 8959
rect 9674 8956 9680 8968
rect 9631 8928 9680 8956
rect 9631 8925 9643 8928
rect 9585 8919 9643 8925
rect 9674 8916 9680 8928
rect 9732 8916 9738 8968
rect 9766 8916 9772 8968
rect 9824 8916 9830 8968
rect 10796 8965 10824 8996
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 11756 8996 12173 9024
rect 11756 8984 11762 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 12434 8984 12440 9036
rect 12492 8984 12498 9036
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 10781 8959 10839 8965
rect 10781 8925 10793 8959
rect 10827 8925 10839 8959
rect 10781 8919 10839 8925
rect 10870 8916 10876 8968
rect 10928 8956 10934 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 10928 8928 11621 8956
rect 10928 8916 10934 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11882 8916 11888 8968
rect 11940 8916 11946 8968
rect 13924 8956 13952 8987
rect 15102 8984 15108 9036
rect 15160 8984 15166 9036
rect 14182 8956 14188 8968
rect 13924 8928 14188 8956
rect 14182 8916 14188 8928
rect 14240 8956 14246 8968
rect 14277 8959 14335 8965
rect 14277 8956 14289 8959
rect 14240 8928 14289 8956
rect 14240 8916 14246 8928
rect 14277 8925 14289 8928
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14366 8916 14372 8968
rect 14424 8916 14430 8968
rect 14642 8916 14648 8968
rect 14700 8916 14706 8968
rect 15120 8941 15148 8984
rect 15105 8935 15163 8941
rect 15105 8901 15117 8935
rect 15151 8901 15163 8935
rect 6181 8891 6239 8897
rect 6181 8857 6193 8891
rect 6227 8888 6239 8891
rect 6549 8891 6607 8897
rect 6549 8888 6561 8891
rect 6227 8860 6561 8888
rect 6227 8857 6239 8860
rect 6181 8851 6239 8857
rect 6549 8857 6561 8860
rect 6595 8857 6607 8891
rect 6549 8851 6607 8857
rect 7558 8848 7564 8900
rect 7616 8848 7622 8900
rect 11333 8891 11391 8897
rect 11333 8857 11345 8891
rect 11379 8857 11391 8891
rect 11333 8851 11391 8857
rect 6638 8820 6644 8832
rect 5920 8792 6644 8820
rect 6638 8780 6644 8792
rect 6696 8820 6702 8832
rect 8021 8823 8079 8829
rect 8021 8820 8033 8823
rect 6696 8792 8033 8820
rect 6696 8780 6702 8792
rect 8021 8789 8033 8792
rect 8067 8789 8079 8823
rect 11348 8820 11376 8851
rect 11422 8848 11428 8900
rect 11480 8888 11486 8900
rect 11701 8891 11759 8897
rect 11701 8888 11713 8891
rect 11480 8860 11713 8888
rect 11480 8848 11486 8860
rect 11701 8857 11713 8860
rect 11747 8888 11759 8891
rect 12342 8888 12348 8900
rect 11747 8860 12348 8888
rect 11747 8857 11759 8860
rect 11701 8851 11759 8857
rect 12342 8848 12348 8860
rect 12400 8848 12406 8900
rect 13170 8848 13176 8900
rect 13228 8848 13234 8900
rect 14458 8848 14464 8900
rect 14516 8848 14522 8900
rect 15105 8895 15163 8901
rect 12158 8820 12164 8832
rect 11348 8792 12164 8820
rect 8021 8783 8079 8789
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 13998 8780 14004 8832
rect 14056 8820 14062 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 14056 8792 14105 8820
rect 14056 8780 14062 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 1104 8730 15456 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 15456 8730
rect 1104 8656 15456 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2314 8616 2320 8628
rect 1811 8588 2320 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2682 8576 2688 8628
rect 2740 8616 2746 8628
rect 4065 8619 4123 8625
rect 4065 8616 4077 8619
rect 2740 8588 4077 8616
rect 2740 8576 2746 8588
rect 4065 8585 4077 8588
rect 4111 8585 4123 8619
rect 4065 8579 4123 8585
rect 4614 8576 4620 8628
rect 4672 8616 4678 8628
rect 4801 8619 4859 8625
rect 4801 8616 4813 8619
rect 4672 8588 4813 8616
rect 4672 8576 4678 8588
rect 4801 8585 4813 8588
rect 4847 8585 4859 8619
rect 4801 8579 4859 8585
rect 4969 8619 5027 8625
rect 4969 8585 4981 8619
rect 5015 8616 5027 8619
rect 5258 8616 5264 8628
rect 5015 8588 5264 8616
rect 5015 8585 5027 8588
rect 4969 8579 5027 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 6546 8616 6552 8628
rect 5776 8588 6552 8616
rect 5776 8576 5782 8588
rect 2130 8508 2136 8560
rect 2188 8548 2194 8560
rect 2225 8551 2283 8557
rect 2225 8548 2237 8551
rect 2188 8520 2237 8548
rect 2188 8508 2194 8520
rect 2225 8517 2237 8520
rect 2271 8517 2283 8551
rect 2225 8511 2283 8517
rect 2869 8551 2927 8557
rect 2869 8517 2881 8551
rect 2915 8548 2927 8551
rect 3050 8548 3056 8560
rect 2915 8520 3056 8548
rect 2915 8517 2927 8520
rect 2869 8511 2927 8517
rect 3050 8508 3056 8520
rect 3108 8508 3114 8560
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 1394 8440 1400 8492
rect 1452 8440 1458 8492
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 4522 8480 4528 8492
rect 2004 8452 4528 8480
rect 2004 8440 2010 8452
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 5074 8440 5080 8492
rect 5132 8480 5138 8492
rect 5184 8480 5212 8511
rect 5350 8508 5356 8560
rect 5408 8548 5414 8560
rect 6472 8557 6500 8588
rect 6546 8576 6552 8588
rect 6604 8576 6610 8628
rect 7098 8576 7104 8628
rect 7156 8576 7162 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7558 8616 7564 8628
rect 7515 8588 7564 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 11330 8576 11336 8628
rect 11388 8576 11394 8628
rect 11514 8576 11520 8628
rect 11572 8616 11578 8628
rect 11675 8619 11733 8625
rect 11675 8616 11687 8619
rect 11572 8588 11687 8616
rect 11572 8576 11578 8588
rect 11675 8585 11687 8588
rect 11721 8585 11733 8619
rect 11675 8579 11733 8585
rect 13814 8576 13820 8628
rect 13872 8576 13878 8628
rect 14461 8619 14519 8625
rect 14461 8585 14473 8619
rect 14507 8616 14519 8619
rect 14642 8616 14648 8628
rect 14507 8588 14648 8616
rect 14507 8585 14519 8588
rect 14461 8579 14519 8585
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 14921 8619 14979 8625
rect 14921 8585 14933 8619
rect 14967 8585 14979 8619
rect 14921 8579 14979 8585
rect 6457 8551 6515 8557
rect 5408 8520 6408 8548
rect 5408 8508 5414 8520
rect 5442 8480 5448 8492
rect 5132 8452 5448 8480
rect 5132 8440 5138 8452
rect 5442 8440 5448 8452
rect 5500 8480 5506 8492
rect 5810 8480 5816 8492
rect 5500 8452 5816 8480
rect 5500 8440 5506 8452
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6380 8489 6408 8520
rect 6457 8517 6469 8551
rect 6503 8548 6515 8551
rect 6503 8520 7328 8548
rect 6503 8517 6515 8520
rect 6457 8511 6515 8517
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8480 6607 8483
rect 6638 8480 6644 8492
rect 6595 8452 6644 8480
rect 6595 8449 6607 8452
rect 6549 8443 6607 8449
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 3016 8415 3074 8421
rect 3016 8412 3028 8415
rect 2832 8384 3028 8412
rect 2832 8372 2838 8384
rect 3016 8381 3028 8384
rect 3062 8381 3074 8415
rect 3016 8375 3074 8381
rect 3237 8415 3295 8421
rect 3237 8381 3249 8415
rect 3283 8412 3295 8415
rect 3326 8412 3332 8424
rect 3283 8384 3332 8412
rect 3283 8381 3295 8384
rect 3237 8375 3295 8381
rect 3326 8372 3332 8384
rect 3384 8372 3390 8424
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3651 8384 3709 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 3973 8415 4031 8421
rect 3973 8412 3985 8415
rect 3936 8384 3985 8412
rect 3936 8372 3942 8384
rect 3973 8381 3985 8384
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 4182 8415 4240 8421
rect 4182 8381 4194 8415
rect 4228 8412 4240 8415
rect 4614 8412 4620 8424
rect 4228 8384 4620 8412
rect 4228 8381 4240 8384
rect 4182 8375 4240 8381
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 5920 8412 5948 8443
rect 6638 8440 6644 8452
rect 6696 8440 6702 8492
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7300 8489 7328 8520
rect 8478 8508 8484 8560
rect 8536 8508 8542 8560
rect 10594 8508 10600 8560
rect 10652 8508 10658 8560
rect 11885 8551 11943 8557
rect 11885 8517 11897 8551
rect 11931 8548 11943 8551
rect 12158 8548 12164 8560
rect 11931 8520 12164 8548
rect 11931 8517 11943 8520
rect 11885 8511 11943 8517
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 13446 8508 13452 8560
rect 13504 8508 13510 8560
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6972 8452 7113 8480
rect 6972 8440 6978 8452
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 7742 8440 7748 8492
rect 7800 8440 7806 8492
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 6454 8412 6460 8424
rect 5920 8384 6460 8412
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 8036 8412 8064 8443
rect 13262 8440 13268 8492
rect 13320 8480 13326 8492
rect 13630 8480 13636 8492
rect 13320 8452 13636 8480
rect 13320 8440 13326 8452
rect 13630 8440 13636 8452
rect 13688 8480 13694 8492
rect 13725 8483 13783 8489
rect 13725 8480 13737 8483
rect 13688 8452 13737 8480
rect 13688 8440 13694 8452
rect 13725 8449 13737 8452
rect 13771 8449 13783 8483
rect 13725 8443 13783 8449
rect 13998 8440 14004 8492
rect 14056 8440 14062 8492
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14274 8440 14280 8492
rect 14332 8440 14338 8492
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8480 14611 8483
rect 14734 8480 14740 8492
rect 14599 8452 14740 8480
rect 14599 8449 14611 8452
rect 14553 8443 14611 8449
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8480 14887 8483
rect 14936 8480 14964 8579
rect 14875 8452 14964 8480
rect 14875 8449 14887 8452
rect 14829 8443 14887 8449
rect 15102 8440 15108 8492
rect 15160 8440 15166 8492
rect 7760 8384 8064 8412
rect 1854 8304 1860 8356
rect 1912 8304 1918 8356
rect 2866 8304 2872 8356
rect 2924 8344 2930 8356
rect 3145 8347 3203 8353
rect 3145 8344 3157 8347
rect 2924 8316 3157 8344
rect 2924 8304 2930 8316
rect 3145 8313 3157 8316
rect 3191 8313 3203 8347
rect 3145 8307 3203 8313
rect 4341 8347 4399 8353
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 7760 8344 7788 8384
rect 9582 8372 9588 8424
rect 9640 8372 9646 8424
rect 9861 8415 9919 8421
rect 9861 8381 9873 8415
rect 9907 8412 9919 8415
rect 9907 8384 11560 8412
rect 9907 8381 9919 8384
rect 9861 8375 9919 8381
rect 11532 8353 11560 8384
rect 4387 8316 7788 8344
rect 7837 8347 7895 8353
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 7837 8313 7849 8347
rect 7883 8313 7895 8347
rect 7837 8307 7895 8313
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8313 11575 8347
rect 11517 8307 11575 8313
rect 1581 8279 1639 8285
rect 1581 8245 1593 8279
rect 1627 8276 1639 8279
rect 1670 8276 1676 8288
rect 1627 8248 1676 8276
rect 1627 8245 1639 8248
rect 1581 8239 1639 8245
rect 1670 8236 1676 8248
rect 1728 8236 1734 8288
rect 4982 8236 4988 8288
rect 5040 8236 5046 8288
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 7852 8276 7880 8307
rect 6328 8248 7880 8276
rect 6328 8236 6334 8248
rect 11422 8236 11428 8288
rect 11480 8276 11486 8288
rect 11701 8279 11759 8285
rect 11701 8276 11713 8279
rect 11480 8248 11713 8276
rect 11480 8236 11486 8248
rect 11701 8245 11713 8248
rect 11747 8245 11759 8279
rect 11701 8239 11759 8245
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 14737 8279 14795 8285
rect 14737 8276 14749 8279
rect 11848 8248 14749 8276
rect 11848 8236 11854 8248
rect 14737 8245 14749 8248
rect 14783 8245 14795 8279
rect 14737 8239 14795 8245
rect 1104 8186 15456 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 15456 8186
rect 1104 8112 15456 8134
rect 4157 8075 4215 8081
rect 4157 8041 4169 8075
rect 4203 8072 4215 8075
rect 4706 8072 4712 8084
rect 4203 8044 4712 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 4706 8032 4712 8044
rect 4764 8032 4770 8084
rect 5074 8032 5080 8084
rect 5132 8032 5138 8084
rect 5261 8075 5319 8081
rect 5261 8041 5273 8075
rect 5307 8072 5319 8075
rect 5350 8072 5356 8084
rect 5307 8044 5356 8072
rect 5307 8041 5319 8044
rect 5261 8035 5319 8041
rect 5350 8032 5356 8044
rect 5408 8032 5414 8084
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 5721 8075 5779 8081
rect 5721 8072 5733 8075
rect 5684 8044 5733 8072
rect 5684 8032 5690 8044
rect 5721 8041 5733 8044
rect 5767 8072 5779 8075
rect 5902 8072 5908 8084
rect 5767 8044 5908 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 7653 8075 7711 8081
rect 7653 8041 7665 8075
rect 7699 8072 7711 8075
rect 7742 8072 7748 8084
rect 7699 8044 7748 8072
rect 7699 8041 7711 8044
rect 7653 8035 7711 8041
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9585 8075 9643 8081
rect 8812 8044 9536 8072
rect 8812 8032 8818 8044
rect 3053 8007 3111 8013
rect 3053 7973 3065 8007
rect 3099 8004 3111 8007
rect 3234 8004 3240 8016
rect 3099 7976 3240 8004
rect 3099 7973 3111 7976
rect 3053 7967 3111 7973
rect 3234 7964 3240 7976
rect 3292 7964 3298 8016
rect 4341 8007 4399 8013
rect 4341 7973 4353 8007
rect 4387 8004 4399 8007
rect 9398 8004 9404 8016
rect 4387 7976 9404 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 4798 7936 4804 7948
rect 2746 7908 4804 7936
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 1946 7828 1952 7880
rect 2004 7828 2010 7880
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2746 7868 2774 7908
rect 4798 7896 4804 7908
rect 4856 7936 4862 7948
rect 4856 7908 4936 7936
rect 4856 7896 4862 7908
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 2280 7840 2774 7868
rect 2976 7840 3341 7868
rect 2280 7828 2286 7840
rect 2038 7760 2044 7812
rect 2096 7800 2102 7812
rect 2682 7800 2688 7812
rect 2096 7772 2688 7800
rect 2096 7760 2102 7772
rect 2682 7760 2688 7772
rect 2740 7800 2746 7812
rect 2976 7800 3004 7840
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3752 7840 3801 7868
rect 3752 7828 3758 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 4908 7809 4936 7908
rect 5350 7896 5356 7948
rect 5408 7896 5414 7948
rect 8036 7945 8064 7976
rect 9398 7964 9404 7976
rect 9456 7964 9462 8016
rect 9508 8004 9536 8044
rect 9585 8041 9597 8075
rect 9631 8072 9643 8075
rect 9766 8072 9772 8084
rect 9631 8044 9772 8072
rect 9631 8041 9643 8044
rect 9585 8035 9643 8041
rect 9766 8032 9772 8044
rect 9824 8032 9830 8084
rect 9950 8032 9956 8084
rect 10008 8072 10014 8084
rect 10008 8044 10272 8072
rect 10008 8032 10014 8044
rect 9858 8004 9864 8016
rect 9508 7976 9864 8004
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 10244 8004 10272 8044
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10689 8075 10747 8081
rect 10689 8072 10701 8075
rect 10652 8044 10701 8072
rect 10652 8032 10658 8044
rect 10689 8041 10701 8044
rect 10735 8041 10747 8075
rect 10689 8035 10747 8041
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 11422 8072 11428 8084
rect 11287 8044 11428 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 11422 8032 11428 8044
rect 11480 8032 11486 8084
rect 14274 8032 14280 8084
rect 14332 8072 14338 8084
rect 14645 8075 14703 8081
rect 14645 8072 14657 8075
rect 14332 8044 14657 8072
rect 14332 8032 14338 8044
rect 14645 8041 14657 8044
rect 14691 8041 14703 8075
rect 14645 8035 14703 8041
rect 14734 8032 14740 8084
rect 14792 8072 14798 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 14792 8044 14933 8072
rect 14792 8032 14798 8044
rect 14921 8041 14933 8044
rect 14967 8041 14979 8075
rect 14921 8035 14979 8041
rect 11790 8004 11796 8016
rect 10244 7976 11796 8004
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 14458 8004 14464 8016
rect 14108 7976 14464 8004
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7905 8079 7939
rect 8021 7899 8079 7905
rect 8665 7939 8723 7945
rect 8665 7905 8677 7939
rect 8711 7936 8723 7939
rect 13354 7936 13360 7948
rect 8711 7908 10088 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7868 7895 7871
rect 7926 7868 7932 7880
rect 7883 7840 7932 7868
rect 7883 7837 7895 7840
rect 7837 7831 7895 7837
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 8754 7828 8760 7880
rect 8812 7828 8818 7880
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7868 8999 7871
rect 8987 7840 9720 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 2740 7772 3004 7800
rect 4893 7803 4951 7809
rect 2740 7760 2746 7772
rect 4893 7769 4905 7803
rect 4939 7769 4951 7803
rect 4893 7763 4951 7769
rect 4982 7760 4988 7812
rect 5040 7800 5046 7812
rect 5093 7803 5151 7809
rect 5093 7800 5105 7803
rect 5040 7772 5105 7800
rect 5040 7760 5046 7772
rect 5093 7769 5105 7772
rect 5139 7800 5151 7803
rect 5258 7800 5264 7812
rect 5139 7772 5264 7800
rect 5139 7769 5151 7772
rect 5093 7763 5151 7769
rect 5258 7760 5264 7772
rect 5316 7760 5322 7812
rect 8297 7803 8355 7809
rect 8297 7769 8309 7803
rect 8343 7800 8355 7803
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8343 7772 9321 7800
rect 8343 7769 8355 7772
rect 8297 7763 8355 7769
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 9398 7760 9404 7812
rect 9456 7809 9462 7812
rect 9456 7803 9484 7809
rect 9472 7769 9484 7803
rect 9456 7763 9484 7769
rect 9456 7760 9462 7763
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 1854 7692 1860 7744
rect 1912 7692 1918 7744
rect 2130 7692 2136 7744
rect 2188 7692 2194 7744
rect 3234 7692 3240 7744
rect 3292 7692 3298 7744
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 3510 7732 3516 7744
rect 3467 7704 3516 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 3510 7692 3516 7704
rect 3568 7692 3574 7744
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 4157 7735 4215 7741
rect 4157 7732 4169 7735
rect 3651 7704 4169 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 4157 7701 4169 7704
rect 4203 7701 4215 7735
rect 4157 7695 4215 7701
rect 5718 7692 5724 7744
rect 5776 7692 5782 7744
rect 5905 7735 5963 7741
rect 5905 7701 5917 7735
rect 5951 7732 5963 7735
rect 7834 7732 7840 7744
rect 5951 7704 7840 7732
rect 5951 7701 5963 7704
rect 5905 7695 5963 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 9122 7692 9128 7744
rect 9180 7732 9186 7744
rect 9692 7741 9720 7840
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 9861 7871 9919 7877
rect 9861 7868 9873 7871
rect 9824 7840 9873 7868
rect 9824 7828 9830 7840
rect 9861 7837 9873 7840
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 10060 7868 10088 7908
rect 10520 7908 13360 7936
rect 10209 7871 10267 7877
rect 10209 7868 10221 7871
rect 10060 7840 10221 7868
rect 10209 7837 10221 7840
rect 10255 7868 10267 7871
rect 10520 7868 10548 7908
rect 13354 7896 13360 7908
rect 13412 7896 13418 7948
rect 10255 7840 10548 7868
rect 10597 7871 10655 7877
rect 10255 7837 10267 7840
rect 10209 7831 10267 7837
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 11057 7871 11115 7877
rect 10643 7840 11008 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 10045 7803 10103 7809
rect 10045 7769 10057 7803
rect 10091 7769 10103 7803
rect 10045 7763 10103 7769
rect 9217 7735 9275 7741
rect 9217 7732 9229 7735
rect 9180 7704 9229 7732
rect 9180 7692 9186 7704
rect 9217 7701 9229 7704
rect 9263 7701 9275 7735
rect 9217 7695 9275 7701
rect 9677 7735 9735 7741
rect 9677 7701 9689 7735
rect 9723 7701 9735 7735
rect 9677 7695 9735 7701
rect 9858 7692 9864 7744
rect 9916 7732 9922 7744
rect 10060 7732 10088 7763
rect 10870 7760 10876 7812
rect 10928 7760 10934 7812
rect 10980 7800 11008 7840
rect 11057 7837 11069 7871
rect 11103 7868 11115 7871
rect 11330 7868 11336 7880
rect 11103 7840 11336 7868
rect 11103 7837 11115 7840
rect 11057 7831 11115 7837
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 14108 7877 14136 7976
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 14185 7939 14243 7945
rect 14185 7905 14197 7939
rect 14231 7936 14243 7939
rect 14642 7936 14648 7948
rect 14231 7908 14648 7936
rect 14231 7905 14243 7908
rect 14185 7899 14243 7905
rect 14642 7896 14648 7908
rect 14700 7896 14706 7948
rect 14093 7871 14151 7877
rect 14093 7837 14105 7871
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7837 14427 7871
rect 14369 7831 14427 7837
rect 11790 7800 11796 7812
rect 10980 7772 11796 7800
rect 11790 7760 11796 7772
rect 11848 7760 11854 7812
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14384 7800 14412 7831
rect 14458 7828 14464 7880
rect 14516 7828 14522 7880
rect 15102 7828 15108 7880
rect 15160 7828 15166 7880
rect 13780 7772 14412 7800
rect 13780 7760 13786 7772
rect 9916 7704 10088 7732
rect 9916 7692 9922 7704
rect 1104 7642 15456 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 15456 7642
rect 1104 7568 15456 7590
rect 2038 7488 2044 7540
rect 2096 7488 2102 7540
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7497 3111 7531
rect 3053 7491 3111 7497
rect 2130 7460 2136 7472
rect 1504 7432 2136 7460
rect 1504 7401 1532 7432
rect 2130 7420 2136 7432
rect 2188 7420 2194 7472
rect 1489 7395 1547 7401
rect 1489 7361 1501 7395
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 1765 7395 1823 7401
rect 1765 7392 1777 7395
rect 1636 7364 1777 7392
rect 1636 7352 1642 7364
rect 1765 7361 1777 7364
rect 1811 7361 1823 7395
rect 1765 7355 1823 7361
rect 1854 7352 1860 7404
rect 1912 7352 1918 7404
rect 2682 7352 2688 7404
rect 2740 7352 2746 7404
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3068 7392 3096 7491
rect 3694 7488 3700 7540
rect 3752 7488 3758 7540
rect 5718 7488 5724 7540
rect 5776 7488 5782 7540
rect 6365 7531 6423 7537
rect 6365 7497 6377 7531
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 3786 7420 3792 7472
rect 3844 7420 3850 7472
rect 4798 7420 4804 7472
rect 4856 7460 4862 7472
rect 5537 7463 5595 7469
rect 5537 7460 5549 7463
rect 4856 7432 5549 7460
rect 4856 7420 4862 7432
rect 5537 7429 5549 7432
rect 5583 7460 5595 7463
rect 6380 7460 6408 7491
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8849 7531 8907 7537
rect 8849 7528 8861 7531
rect 7984 7500 8861 7528
rect 7984 7488 7990 7500
rect 8849 7497 8861 7500
rect 8895 7497 8907 7531
rect 8849 7491 8907 7497
rect 9122 7488 9128 7540
rect 9180 7488 9186 7540
rect 5583 7432 6408 7460
rect 5583 7429 5595 7432
rect 5537 7423 5595 7429
rect 7834 7420 7840 7472
rect 7892 7420 7898 7472
rect 8386 7469 8392 7472
rect 8363 7463 8392 7469
rect 8363 7429 8375 7463
rect 8363 7423 8392 7429
rect 8386 7420 8392 7423
rect 8444 7420 8450 7472
rect 9309 7463 9367 7469
rect 9309 7429 9321 7463
rect 9355 7460 9367 7463
rect 9950 7460 9956 7472
rect 9355 7432 9956 7460
rect 9355 7429 9367 7432
rect 9309 7423 9367 7429
rect 9950 7420 9956 7432
rect 10008 7420 10014 7472
rect 13633 7463 13691 7469
rect 13633 7460 13645 7463
rect 13202 7432 13645 7460
rect 13633 7429 13645 7432
rect 13679 7429 13691 7463
rect 13633 7423 13691 7429
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 3068 7364 3341 7392
rect 3329 7361 3341 7364
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7392 3571 7395
rect 3878 7392 3884 7404
rect 3559 7364 3884 7392
rect 3559 7361 3571 7364
rect 3513 7355 3571 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 5350 7352 5356 7404
rect 5408 7352 5414 7404
rect 6730 7352 6736 7404
rect 6788 7352 6794 7404
rect 8478 7352 8484 7404
rect 8536 7352 8542 7404
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 8665 7395 8723 7401
rect 8665 7361 8677 7395
rect 8711 7392 8723 7395
rect 9122 7392 9128 7404
rect 8711 7364 9128 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 2133 7327 2191 7333
rect 2133 7293 2145 7327
rect 2179 7324 2191 7327
rect 2222 7324 2228 7336
rect 2179 7296 2228 7324
rect 2179 7293 2191 7296
rect 2133 7287 2191 7293
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2593 7327 2651 7333
rect 2593 7293 2605 7327
rect 2639 7324 2651 7327
rect 2884 7324 2912 7352
rect 2639 7296 2912 7324
rect 8113 7327 8171 7333
rect 2639 7293 2651 7296
rect 2593 7287 2651 7293
rect 8113 7293 8125 7327
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 1670 7256 1676 7268
rect 1627 7228 1676 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 1670 7216 1676 7228
rect 1728 7256 1734 7268
rect 2409 7259 2467 7265
rect 2409 7256 2421 7259
rect 1728 7228 2421 7256
rect 1728 7216 1734 7228
rect 2409 7225 2421 7228
rect 2455 7225 2467 7259
rect 2409 7219 2467 7225
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3789 7259 3847 7265
rect 3789 7256 3801 7259
rect 3292 7228 3801 7256
rect 3292 7216 3298 7228
rect 3789 7225 3801 7228
rect 3835 7225 3847 7259
rect 3789 7219 3847 7225
rect 2774 7148 2780 7200
rect 2832 7148 2838 7200
rect 3326 7148 3332 7200
rect 3384 7148 3390 7200
rect 8128 7188 8156 7287
rect 8202 7284 8208 7336
rect 8260 7284 8266 7336
rect 8588 7324 8616 7355
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 8846 7324 8852 7336
rect 8588 7296 8852 7324
rect 8846 7284 8852 7296
rect 8904 7284 8910 7336
rect 9508 7256 9536 7355
rect 9582 7352 9588 7404
rect 9640 7392 9646 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9640 7364 10333 7392
rect 9640 7352 9646 7364
rect 10321 7361 10333 7364
rect 10367 7392 10379 7395
rect 11698 7392 11704 7404
rect 10367 7364 11704 7392
rect 10367 7361 10379 7364
rect 10321 7355 10379 7361
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7361 13783 7395
rect 13725 7355 13783 7361
rect 11974 7284 11980 7336
rect 12032 7284 12038 7336
rect 9766 7256 9772 7268
rect 9508 7228 9772 7256
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 13740 7256 13768 7355
rect 14458 7352 14464 7404
rect 14516 7352 14522 7404
rect 14737 7395 14795 7401
rect 14737 7392 14749 7395
rect 14660 7364 14749 7392
rect 14660 7265 14688 7364
rect 14737 7361 14749 7364
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 13096 7228 13768 7256
rect 14645 7259 14703 7265
rect 9582 7188 9588 7200
rect 8128 7160 9588 7188
rect 9582 7148 9588 7160
rect 9640 7148 9646 7200
rect 11790 7148 11796 7200
rect 11848 7188 11854 7200
rect 13096 7188 13124 7228
rect 14645 7225 14657 7259
rect 14691 7225 14703 7259
rect 14645 7219 14703 7225
rect 11848 7160 13124 7188
rect 11848 7148 11854 7160
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13449 7191 13507 7197
rect 13449 7188 13461 7191
rect 13228 7160 13461 7188
rect 13228 7148 13234 7160
rect 13449 7157 13461 7160
rect 13495 7188 13507 7191
rect 13722 7188 13728 7200
rect 13495 7160 13728 7188
rect 13495 7157 13507 7160
rect 13449 7151 13507 7157
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 14829 7191 14887 7197
rect 14829 7188 14841 7191
rect 14424 7160 14841 7188
rect 14424 7148 14430 7160
rect 14829 7157 14841 7160
rect 14875 7157 14887 7191
rect 14829 7151 14887 7157
rect 1104 7098 15456 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 15456 7098
rect 1104 7024 15456 7046
rect 3881 6987 3939 6993
rect 3881 6953 3893 6987
rect 3927 6984 3939 6987
rect 3970 6984 3976 6996
rect 3927 6956 3976 6984
rect 3927 6953 3939 6956
rect 3881 6947 3939 6953
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 5350 6944 5356 6996
rect 5408 6984 5414 6996
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 5408 6956 5457 6984
rect 5408 6944 5414 6956
rect 5445 6953 5457 6956
rect 5491 6953 5503 6987
rect 5445 6947 5503 6953
rect 5721 6987 5779 6993
rect 5721 6953 5733 6987
rect 5767 6984 5779 6987
rect 5994 6984 6000 6996
rect 5767 6956 6000 6984
rect 5767 6953 5779 6956
rect 5721 6947 5779 6953
rect 5994 6944 6000 6956
rect 6052 6944 6058 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8389 6987 8447 6993
rect 8389 6984 8401 6987
rect 8352 6956 8401 6984
rect 8352 6944 8358 6956
rect 8389 6953 8401 6956
rect 8435 6953 8447 6987
rect 8389 6947 8447 6953
rect 8478 6944 8484 6996
rect 8536 6984 8542 6996
rect 8573 6987 8631 6993
rect 8573 6984 8585 6987
rect 8536 6956 8585 6984
rect 8536 6944 8542 6956
rect 8573 6953 8585 6956
rect 8619 6953 8631 6987
rect 8573 6947 8631 6953
rect 11698 6944 11704 6996
rect 11756 6944 11762 6996
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 12032 6956 12081 6984
rect 12032 6944 12038 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 12216 6956 12265 6984
rect 12216 6944 12222 6956
rect 12253 6953 12265 6956
rect 12299 6953 12311 6987
rect 12253 6947 12311 6953
rect 1578 6876 1584 6928
rect 1636 6916 1642 6928
rect 2041 6919 2099 6925
rect 2041 6916 2053 6919
rect 1636 6888 2053 6916
rect 1636 6876 1642 6888
rect 2041 6885 2053 6888
rect 2087 6885 2099 6919
rect 8021 6919 8079 6925
rect 2041 6879 2099 6885
rect 6656 6888 7052 6916
rect 1765 6851 1823 6857
rect 1765 6817 1777 6851
rect 1811 6848 1823 6851
rect 1946 6848 1952 6860
rect 1811 6820 1952 6848
rect 1811 6817 1823 6820
rect 1765 6811 1823 6817
rect 1946 6808 1952 6820
rect 2004 6808 2010 6860
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2774 6848 2780 6860
rect 2271 6820 2780 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 5077 6851 5135 6857
rect 5077 6817 5089 6851
rect 5123 6848 5135 6851
rect 5442 6848 5448 6860
rect 5123 6820 5448 6848
rect 5123 6817 5135 6820
rect 5077 6811 5135 6817
rect 5442 6808 5448 6820
rect 5500 6848 5506 6860
rect 6656 6848 6684 6888
rect 5500 6820 6684 6848
rect 5500 6808 5506 6820
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 6917 6851 6975 6857
rect 6917 6848 6929 6851
rect 6788 6820 6929 6848
rect 6788 6808 6794 6820
rect 6917 6817 6929 6820
rect 6963 6817 6975 6851
rect 7024 6848 7052 6888
rect 8021 6885 8033 6919
rect 8067 6916 8079 6919
rect 8202 6916 8208 6928
rect 8067 6888 8208 6916
rect 8067 6885 8079 6888
rect 8021 6879 8079 6885
rect 8202 6876 8208 6888
rect 8260 6876 8266 6928
rect 10870 6876 10876 6928
rect 10928 6916 10934 6928
rect 10928 6888 12434 6916
rect 10928 6876 10934 6888
rect 7024 6820 7696 6848
rect 6917 6811 6975 6817
rect 3973 6783 4031 6789
rect 3973 6749 3985 6783
rect 4019 6780 4031 6783
rect 4246 6780 4252 6792
rect 4019 6752 4252 6780
rect 4019 6749 4031 6752
rect 3973 6743 4031 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6780 6883 6783
rect 7558 6780 7564 6792
rect 6871 6752 7564 6780
rect 6871 6749 6883 6752
rect 6825 6743 6883 6749
rect 5276 6644 5304 6740
rect 6932 6724 6960 6752
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7668 6780 7696 6820
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9306 6848 9312 6860
rect 8812 6820 9312 6848
rect 8812 6808 8818 6820
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 12406 6848 12434 6888
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12406 6820 12633 6848
rect 12621 6817 12633 6820
rect 12667 6848 12679 6851
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 12667 6820 13369 6848
rect 12667 6817 12679 6820
rect 12621 6811 12679 6817
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 9122 6780 9128 6792
rect 7668 6752 9128 6780
rect 9122 6740 9128 6752
rect 9180 6780 9186 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9180 6752 9505 6780
rect 9180 6740 9186 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12768 6752 12909 6780
rect 12768 6740 12774 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 12986 6740 12992 6792
rect 13044 6740 13050 6792
rect 13081 6783 13139 6789
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 5905 6715 5963 6721
rect 5905 6681 5917 6715
rect 5951 6712 5963 6715
rect 6086 6712 6092 6724
rect 5951 6684 6092 6712
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 6914 6672 6920 6724
rect 6972 6672 6978 6724
rect 8938 6672 8944 6724
rect 8996 6712 9002 6724
rect 10229 6715 10287 6721
rect 10229 6712 10241 6715
rect 8996 6684 10241 6712
rect 8996 6672 9002 6684
rect 10229 6681 10241 6684
rect 10275 6681 10287 6715
rect 10229 6675 10287 6681
rect 12434 6672 12440 6724
rect 12492 6712 12498 6724
rect 13096 6712 13124 6743
rect 13170 6740 13176 6792
rect 13228 6740 13234 6792
rect 13538 6740 13544 6792
rect 13596 6740 13602 6792
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 13909 6783 13967 6789
rect 13909 6780 13921 6783
rect 13780 6752 13921 6780
rect 13780 6740 13786 6752
rect 13909 6749 13921 6752
rect 13955 6780 13967 6783
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 13955 6752 14289 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14366 6740 14372 6792
rect 14424 6740 14430 6792
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 14461 6715 14519 6721
rect 12492 6684 14412 6712
rect 12492 6672 12498 6684
rect 13740 6656 13768 6684
rect 5718 6653 5724 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 5276 6616 5549 6644
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5537 6607 5595 6613
rect 5705 6647 5724 6653
rect 5705 6613 5717 6647
rect 5705 6607 5724 6613
rect 5718 6604 5724 6607
rect 5776 6604 5782 6656
rect 8386 6604 8392 6656
rect 8444 6604 8450 6656
rect 9674 6604 9680 6656
rect 9732 6604 9738 6656
rect 12253 6647 12311 6653
rect 12253 6613 12265 6647
rect 12299 6644 12311 6647
rect 12713 6647 12771 6653
rect 12713 6644 12725 6647
rect 12299 6616 12725 6644
rect 12299 6613 12311 6616
rect 12253 6607 12311 6613
rect 12713 6613 12725 6616
rect 12759 6613 12771 6647
rect 12713 6607 12771 6613
rect 12986 6604 12992 6656
rect 13044 6644 13050 6656
rect 13446 6644 13452 6656
rect 13044 6616 13452 6644
rect 13044 6604 13050 6616
rect 13446 6604 13452 6616
rect 13504 6604 13510 6656
rect 13630 6604 13636 6656
rect 13688 6604 13694 6656
rect 13722 6604 13728 6656
rect 13780 6604 13786 6656
rect 14090 6604 14096 6656
rect 14148 6604 14154 6656
rect 14384 6644 14412 6684
rect 14461 6681 14473 6715
rect 14507 6712 14519 6715
rect 14550 6712 14556 6724
rect 14507 6684 14556 6712
rect 14507 6681 14519 6684
rect 14461 6675 14519 6681
rect 14550 6672 14556 6684
rect 14608 6672 14614 6724
rect 14660 6644 14688 6743
rect 15102 6740 15108 6792
rect 15160 6740 15166 6792
rect 14384 6616 14688 6644
rect 14918 6604 14924 6656
rect 14976 6604 14982 6656
rect 1104 6554 15456 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 15456 6554
rect 1104 6480 15456 6502
rect 2501 6443 2559 6449
rect 2501 6409 2513 6443
rect 2547 6440 2559 6443
rect 2682 6440 2688 6452
rect 2547 6412 2688 6440
rect 2547 6409 2559 6412
rect 2501 6403 2559 6409
rect 2682 6400 2688 6412
rect 2740 6440 2746 6452
rect 3237 6443 3295 6449
rect 2740 6400 2774 6440
rect 3237 6409 3249 6443
rect 3283 6440 3295 6443
rect 4614 6440 4620 6452
rect 3283 6412 4620 6440
rect 3283 6409 3295 6412
rect 3237 6403 3295 6409
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 8202 6400 8208 6452
rect 8260 6400 8266 6452
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 9364 6412 9597 6440
rect 9364 6400 9370 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 11609 6443 11667 6449
rect 11609 6409 11621 6443
rect 11655 6409 11667 6443
rect 11609 6403 11667 6409
rect 13449 6443 13507 6449
rect 13449 6409 13461 6443
rect 13495 6440 13507 6443
rect 14182 6440 14188 6452
rect 13495 6412 14188 6440
rect 13495 6409 13507 6412
rect 13449 6403 13507 6409
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 2593 6307 2651 6313
rect 2593 6304 2605 6307
rect 1397 6267 1455 6273
rect 1964 6276 2605 6304
rect 1581 6171 1639 6177
rect 1581 6137 1593 6171
rect 1627 6168 1639 6171
rect 1964 6168 1992 6276
rect 2593 6273 2605 6276
rect 2639 6273 2651 6307
rect 2746 6304 2774 6400
rect 3973 6375 4031 6381
rect 3973 6341 3985 6375
rect 4019 6372 4031 6375
rect 4062 6372 4068 6384
rect 4019 6344 4068 6372
rect 4019 6341 4031 6344
rect 3973 6335 4031 6341
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 5626 6332 5632 6384
rect 5684 6332 5690 6384
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 9324 6372 9352 6400
rect 11624 6372 11652 6403
rect 14182 6400 14188 6412
rect 14240 6400 14246 6452
rect 9088 6344 9352 6372
rect 10626 6344 11652 6372
rect 12345 6375 12403 6381
rect 9088 6332 9094 6344
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 2746 6276 3433 6304
rect 2593 6267 2651 6273
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3510 6264 3516 6316
rect 3568 6304 3574 6316
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3568 6276 3709 6304
rect 3568 6264 3574 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6304 3939 6307
rect 4525 6307 4583 6313
rect 4525 6304 4537 6307
rect 3927 6276 4537 6304
rect 3927 6273 3939 6276
rect 3881 6267 3939 6273
rect 4525 6273 4537 6276
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 2041 6239 2099 6245
rect 2041 6205 2053 6239
rect 2087 6236 2099 6239
rect 4724 6236 4752 6267
rect 4890 6264 4896 6316
rect 4948 6264 4954 6316
rect 4982 6264 4988 6316
rect 5040 6264 5046 6316
rect 5261 6307 5319 6313
rect 5261 6273 5273 6307
rect 5307 6304 5319 6307
rect 5350 6304 5356 6316
rect 5307 6276 5356 6304
rect 5307 6273 5319 6276
rect 5261 6267 5319 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 6730 6264 6736 6316
rect 6788 6264 6794 6316
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8481 6307 8539 6313
rect 8481 6304 8493 6307
rect 8260 6276 8493 6304
rect 8260 6264 8266 6276
rect 8481 6273 8493 6276
rect 8527 6273 8539 6307
rect 8481 6267 8539 6273
rect 9122 6264 9128 6316
rect 9180 6264 9186 6316
rect 9324 6313 9352 6344
rect 12345 6341 12357 6375
rect 12391 6372 12403 6375
rect 12986 6372 12992 6384
rect 12391 6344 12992 6372
rect 12391 6341 12403 6344
rect 12345 6335 12403 6341
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 14090 6372 14096 6384
rect 13648 6344 14096 6372
rect 9309 6307 9367 6313
rect 9309 6273 9321 6307
rect 9355 6273 9367 6307
rect 9309 6267 9367 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11606 6304 11612 6316
rect 11379 6276 11612 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 11790 6304 11796 6316
rect 11747 6276 11796 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 12161 6307 12219 6313
rect 12161 6273 12173 6307
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 7837 6239 7895 6245
rect 7837 6236 7849 6239
rect 2087 6208 2544 6236
rect 2087 6205 2099 6208
rect 2041 6199 2099 6205
rect 2317 6171 2375 6177
rect 2317 6168 2329 6171
rect 1627 6140 2329 6168
rect 1627 6137 1639 6140
rect 1581 6131 1639 6137
rect 2317 6137 2329 6140
rect 2363 6137 2375 6171
rect 2516 6168 2544 6208
rect 4172 6208 4752 6236
rect 5828 6208 7849 6236
rect 2866 6168 2872 6180
rect 2516 6140 2872 6168
rect 2317 6131 2375 6137
rect 2866 6128 2872 6140
rect 2924 6128 2930 6180
rect 4172 6168 4200 6208
rect 3068 6140 4200 6168
rect 3068 6112 3096 6140
rect 4246 6128 4252 6180
rect 4304 6128 4310 6180
rect 4433 6171 4491 6177
rect 4433 6137 4445 6171
rect 4479 6168 4491 6171
rect 4614 6168 4620 6180
rect 4479 6140 4620 6168
rect 4479 6137 4491 6140
rect 4433 6131 4491 6137
rect 4614 6128 4620 6140
rect 4672 6128 4678 6180
rect 5828 6177 5856 6208
rect 7837 6205 7849 6208
rect 7883 6205 7895 6239
rect 7837 6199 7895 6205
rect 8113 6239 8171 6245
rect 8113 6205 8125 6239
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8570 6236 8576 6248
rect 8435 6208 8576 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 5813 6171 5871 6177
rect 5813 6137 5825 6171
rect 5859 6137 5871 6171
rect 5813 6131 5871 6137
rect 3050 6060 3056 6112
rect 3108 6060 3114 6112
rect 4264 6100 4292 6128
rect 5258 6100 5264 6112
rect 4264 6072 5264 6100
rect 5258 6060 5264 6072
rect 5316 6060 5322 6112
rect 5629 6103 5687 6109
rect 5629 6069 5641 6103
rect 5675 6100 5687 6103
rect 5902 6100 5908 6112
rect 5675 6072 5908 6100
rect 5675 6069 5687 6072
rect 5629 6063 5687 6069
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6086 6060 6092 6112
rect 6144 6100 6150 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 6144 6072 6377 6100
rect 6144 6060 6150 6072
rect 6365 6069 6377 6072
rect 6411 6069 6423 6103
rect 6365 6063 6423 6069
rect 6822 6060 6828 6112
rect 6880 6100 6886 6112
rect 8128 6100 8156 6199
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 8754 6196 8760 6248
rect 8812 6196 8818 6248
rect 8846 6196 8852 6248
rect 8904 6196 8910 6248
rect 11054 6196 11060 6248
rect 11112 6196 11118 6248
rect 12176 6236 12204 6267
rect 12434 6264 12440 6316
rect 12492 6264 12498 6316
rect 13648 6313 13676 6344
rect 14090 6332 14096 6344
rect 14148 6332 14154 6384
rect 14366 6372 14372 6384
rect 14200 6344 14372 6372
rect 13173 6307 13231 6313
rect 13173 6273 13185 6307
rect 13219 6273 13231 6307
rect 13173 6267 13231 6273
rect 13633 6307 13691 6313
rect 13633 6273 13645 6307
rect 13679 6273 13691 6307
rect 13633 6267 13691 6273
rect 12618 6236 12624 6248
rect 12176 6208 12624 6236
rect 12618 6196 12624 6208
rect 12676 6196 12682 6248
rect 13188 6236 13216 6267
rect 13814 6264 13820 6316
rect 13872 6264 13878 6316
rect 14200 6313 14228 6344
rect 14366 6332 14372 6344
rect 14424 6372 14430 6384
rect 14829 6375 14887 6381
rect 14829 6372 14841 6375
rect 14424 6344 14841 6372
rect 14424 6332 14430 6344
rect 14829 6341 14841 6344
rect 14875 6341 14887 6375
rect 14829 6335 14887 6341
rect 13909 6307 13967 6313
rect 13909 6273 13921 6307
rect 13955 6304 13967 6307
rect 14001 6307 14059 6313
rect 14001 6304 14013 6307
rect 13955 6276 14013 6304
rect 13955 6273 13967 6276
rect 13909 6267 13967 6273
rect 14001 6273 14013 6276
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6273 14243 6307
rect 14185 6267 14243 6273
rect 14274 6264 14280 6316
rect 14332 6264 14338 6316
rect 14550 6264 14556 6316
rect 14608 6264 14614 6316
rect 14918 6264 14924 6316
rect 14976 6264 14982 6316
rect 15194 6236 15200 6248
rect 13188 6208 15200 6236
rect 15194 6196 15200 6208
rect 15252 6196 15258 6248
rect 12158 6168 12164 6180
rect 11900 6140 12164 6168
rect 6880 6072 8156 6100
rect 6880 6060 6886 6072
rect 9490 6060 9496 6112
rect 9548 6060 9554 6112
rect 9950 6060 9956 6112
rect 10008 6100 10014 6112
rect 11900 6100 11928 6140
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 13357 6171 13415 6177
rect 13357 6137 13369 6171
rect 13403 6168 13415 6171
rect 14734 6168 14740 6180
rect 13403 6140 14740 6168
rect 13403 6137 13415 6140
rect 13357 6131 13415 6137
rect 14734 6128 14740 6140
rect 14792 6128 14798 6180
rect 10008 6072 11928 6100
rect 10008 6060 10014 6072
rect 11974 6060 11980 6112
rect 12032 6100 12038 6112
rect 12253 6103 12311 6109
rect 12253 6100 12265 6103
rect 12032 6072 12265 6100
rect 12032 6060 12038 6072
rect 12253 6069 12265 6072
rect 12299 6069 12311 6103
rect 12253 6063 12311 6069
rect 13722 6060 13728 6112
rect 13780 6100 13786 6112
rect 14461 6103 14519 6109
rect 14461 6100 14473 6103
rect 13780 6072 14473 6100
rect 13780 6060 13786 6072
rect 14461 6069 14473 6072
rect 14507 6069 14519 6103
rect 14461 6063 14519 6069
rect 1104 6010 15456 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 15456 6010
rect 1104 5936 15456 5958
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 3878 5896 3884 5908
rect 3835 5868 3884 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4157 5899 4215 5905
rect 4157 5865 4169 5899
rect 4203 5896 4215 5899
rect 4614 5896 4620 5908
rect 4203 5868 4620 5896
rect 4203 5865 4215 5868
rect 4157 5859 4215 5865
rect 4614 5856 4620 5868
rect 4672 5856 4678 5908
rect 5353 5899 5411 5905
rect 5353 5865 5365 5899
rect 5399 5896 5411 5899
rect 5626 5896 5632 5908
rect 5399 5868 5632 5896
rect 5399 5865 5411 5868
rect 5353 5859 5411 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8941 5899 8999 5905
rect 8941 5896 8953 5899
rect 8444 5868 8953 5896
rect 8444 5856 8450 5868
rect 8941 5865 8953 5868
rect 8987 5865 8999 5899
rect 8941 5859 8999 5865
rect 9048 5868 9812 5896
rect 3050 5788 3056 5840
rect 3108 5828 3114 5840
rect 4249 5831 4307 5837
rect 4249 5828 4261 5831
rect 3108 5800 4261 5828
rect 3108 5788 3114 5800
rect 4249 5797 4261 5800
rect 4295 5797 4307 5831
rect 5718 5828 5724 5840
rect 4249 5791 4307 5797
rect 5552 5800 5724 5828
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4706 5760 4712 5772
rect 4111 5732 4712 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4706 5720 4712 5732
rect 4764 5720 4770 5772
rect 5552 5769 5580 5800
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 5902 5788 5908 5840
rect 5960 5828 5966 5840
rect 9048 5828 9076 5868
rect 5960 5800 9076 5828
rect 9585 5831 9643 5837
rect 5960 5788 5966 5800
rect 9585 5797 9597 5831
rect 9631 5828 9643 5831
rect 9674 5828 9680 5840
rect 9631 5800 9680 5828
rect 9631 5797 9643 5800
rect 9585 5791 9643 5797
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 5537 5763 5595 5769
rect 5537 5729 5549 5763
rect 5583 5729 5595 5763
rect 5537 5723 5595 5729
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 5994 5760 6000 5772
rect 5675 5732 6000 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 5994 5720 6000 5732
rect 6052 5720 6058 5772
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4798 5692 4804 5704
rect 4571 5664 4804 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4798 5652 4804 5664
rect 4856 5692 4862 5704
rect 4982 5692 4988 5704
rect 4856 5664 4988 5692
rect 4856 5652 4862 5664
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5442 5652 5448 5704
rect 5500 5692 5506 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5500 5664 5733 5692
rect 5500 5652 5506 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 6086 5692 6092 5704
rect 5859 5664 6092 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 2866 5584 2872 5636
rect 2924 5624 2930 5636
rect 5828 5624 5856 5655
rect 6086 5652 6092 5664
rect 6144 5652 6150 5704
rect 6178 5652 6184 5704
rect 6236 5692 6242 5704
rect 6457 5695 6515 5701
rect 6457 5692 6469 5695
rect 6236 5664 6469 5692
rect 6236 5652 6242 5664
rect 6457 5661 6469 5664
rect 6503 5692 6515 5695
rect 6822 5692 6828 5704
rect 6503 5664 6828 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 6822 5652 6828 5664
rect 6880 5652 6886 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 8938 5692 8944 5704
rect 8619 5664 8944 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9692 5692 9720 5788
rect 9784 5760 9812 5868
rect 9950 5856 9956 5908
rect 10008 5856 10014 5908
rect 10137 5899 10195 5905
rect 10137 5865 10149 5899
rect 10183 5896 10195 5899
rect 11054 5896 11060 5908
rect 10183 5868 11060 5896
rect 10183 5865 10195 5868
rect 10137 5859 10195 5865
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11882 5856 11888 5908
rect 11940 5856 11946 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12526 5896 12532 5908
rect 12124 5868 12532 5896
rect 12124 5856 12130 5868
rect 12526 5856 12532 5868
rect 12584 5856 12590 5908
rect 13814 5856 13820 5908
rect 13872 5896 13878 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13872 5868 14105 5896
rect 13872 5856 13878 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 14550 5856 14556 5908
rect 14608 5896 14614 5908
rect 14829 5899 14887 5905
rect 14829 5896 14841 5899
rect 14608 5868 14841 5896
rect 14608 5856 14614 5868
rect 14829 5865 14841 5868
rect 14875 5865 14887 5899
rect 14829 5859 14887 5865
rect 13722 5788 13728 5840
rect 13780 5828 13786 5840
rect 13909 5831 13967 5837
rect 13909 5828 13921 5831
rect 13780 5800 13921 5828
rect 13780 5788 13786 5800
rect 13909 5797 13921 5800
rect 13955 5797 13967 5831
rect 13909 5791 13967 5797
rect 9784 5732 10364 5760
rect 10229 5695 10287 5701
rect 10229 5692 10241 5695
rect 9692 5664 10241 5692
rect 10229 5661 10241 5664
rect 10275 5661 10287 5695
rect 10336 5692 10364 5732
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 11756 5732 12173 5760
rect 11756 5720 11762 5732
rect 12161 5729 12173 5732
rect 12207 5760 12219 5763
rect 12986 5760 12992 5772
rect 12207 5732 12992 5760
rect 12207 5729 12219 5732
rect 12161 5723 12219 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 12066 5692 12072 5704
rect 10336 5664 12072 5692
rect 10229 5655 10287 5661
rect 2924 5596 5856 5624
rect 2924 5584 2930 5596
rect 8478 5584 8484 5636
rect 8536 5624 8542 5636
rect 8846 5624 8852 5636
rect 8536 5596 8852 5624
rect 8536 5584 8542 5596
rect 8846 5584 8852 5596
rect 8904 5624 8910 5636
rect 9125 5627 9183 5633
rect 9125 5624 9137 5627
rect 8904 5596 9137 5624
rect 8904 5584 8910 5596
rect 9125 5593 9137 5596
rect 9171 5593 9183 5627
rect 9125 5587 9183 5593
rect 9309 5627 9367 5633
rect 9309 5593 9321 5627
rect 9355 5593 9367 5627
rect 9309 5587 9367 5593
rect 4433 5559 4491 5565
rect 4433 5525 4445 5559
rect 4479 5556 4491 5559
rect 4614 5556 4620 5568
rect 4479 5528 4620 5556
rect 4479 5525 4491 5528
rect 4433 5519 4491 5525
rect 4614 5516 4620 5528
rect 4672 5556 4678 5568
rect 4890 5556 4896 5568
rect 4672 5528 4896 5556
rect 4672 5516 4678 5528
rect 4890 5516 4896 5528
rect 4948 5516 4954 5568
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 8938 5556 8944 5568
rect 8812 5528 8944 5556
rect 8812 5516 8818 5528
rect 8938 5516 8944 5528
rect 8996 5556 9002 5568
rect 9324 5556 9352 5587
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 9953 5627 10011 5633
rect 9953 5624 9965 5627
rect 9548 5596 9965 5624
rect 9548 5584 9554 5596
rect 9953 5593 9965 5596
rect 9999 5593 10011 5627
rect 9953 5587 10011 5593
rect 10413 5627 10471 5633
rect 10413 5593 10425 5627
rect 10459 5624 10471 5627
rect 10502 5624 10508 5636
rect 10459 5596 10508 5624
rect 10459 5593 10471 5596
rect 10413 5587 10471 5593
rect 10502 5584 10508 5596
rect 10560 5584 10566 5636
rect 11716 5633 11744 5664
rect 12066 5652 12072 5664
rect 12124 5652 12130 5704
rect 13722 5652 13728 5704
rect 13780 5692 13786 5704
rect 14274 5692 14280 5704
rect 13780 5664 14280 5692
rect 13780 5652 13786 5664
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 14366 5652 14372 5704
rect 14424 5652 14430 5704
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14645 5695 14703 5701
rect 14645 5661 14657 5695
rect 14691 5661 14703 5695
rect 14645 5655 14703 5661
rect 11974 5633 11980 5636
rect 11701 5627 11759 5633
rect 11701 5593 11713 5627
rect 11747 5593 11759 5627
rect 11701 5587 11759 5593
rect 11917 5627 11980 5633
rect 11917 5593 11929 5627
rect 11963 5593 11980 5627
rect 11917 5587 11980 5593
rect 11974 5584 11980 5587
rect 12032 5584 12038 5636
rect 12437 5627 12495 5633
rect 12437 5593 12449 5627
rect 12483 5593 12495 5627
rect 13814 5624 13820 5636
rect 13662 5596 13820 5624
rect 12437 5587 12495 5593
rect 8996 5528 9352 5556
rect 8996 5516 9002 5528
rect 10594 5516 10600 5568
rect 10652 5516 10658 5568
rect 12069 5559 12127 5565
rect 12069 5525 12081 5559
rect 12115 5556 12127 5559
rect 12452 5556 12480 5587
rect 13814 5584 13820 5596
rect 13872 5584 13878 5636
rect 12115 5528 12480 5556
rect 12115 5525 12127 5528
rect 12069 5519 12127 5525
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 13354 5556 13360 5568
rect 12676 5528 13360 5556
rect 12676 5516 12682 5528
rect 13354 5516 13360 5528
rect 13412 5556 13418 5568
rect 14660 5556 14688 5655
rect 14734 5652 14740 5704
rect 14792 5652 14798 5704
rect 13412 5528 14688 5556
rect 13412 5516 13418 5528
rect 1104 5466 15456 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 15456 5466
rect 1104 5392 15456 5414
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 6917 5355 6975 5361
rect 6917 5352 6929 5355
rect 6788 5324 6929 5352
rect 6788 5312 6794 5324
rect 6917 5321 6929 5324
rect 6963 5321 6975 5355
rect 6917 5315 6975 5321
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 8294 5352 8300 5364
rect 8067 5324 8300 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 8849 5355 8907 5361
rect 8849 5321 8861 5355
rect 8895 5352 8907 5355
rect 9030 5352 9036 5364
rect 8895 5324 9036 5352
rect 8895 5321 8907 5324
rect 8849 5315 8907 5321
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9122 5312 9128 5364
rect 9180 5352 9186 5364
rect 9283 5355 9341 5361
rect 9283 5352 9295 5355
rect 9180 5324 9295 5352
rect 9180 5312 9186 5324
rect 9283 5321 9295 5324
rect 9329 5321 9341 5355
rect 9766 5352 9772 5364
rect 9283 5315 9341 5321
rect 9508 5324 9772 5352
rect 8570 5284 8576 5296
rect 8128 5256 8576 5284
rect 8128 5228 8156 5256
rect 8570 5244 8576 5256
rect 8628 5244 8634 5296
rect 8665 5287 8723 5293
rect 8665 5253 8677 5287
rect 8711 5284 8723 5287
rect 8938 5284 8944 5296
rect 8711 5256 8944 5284
rect 8711 5253 8723 5256
rect 8665 5247 8723 5253
rect 8938 5244 8944 5256
rect 8996 5244 9002 5296
rect 9508 5293 9536 5324
rect 9766 5312 9772 5324
rect 9824 5352 9830 5364
rect 10502 5352 10508 5364
rect 9824 5324 10508 5352
rect 9824 5312 9830 5324
rect 10502 5312 10508 5324
rect 10560 5352 10566 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 10560 5324 11345 5352
rect 10560 5312 10566 5324
rect 11333 5321 11345 5324
rect 11379 5321 11391 5355
rect 11333 5315 11391 5321
rect 11882 5312 11888 5364
rect 11940 5352 11946 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11940 5324 12173 5352
rect 11940 5312 11946 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 12529 5355 12587 5361
rect 12529 5321 12541 5355
rect 12575 5352 12587 5355
rect 13722 5352 13728 5364
rect 12575 5324 13728 5352
rect 12575 5321 12587 5324
rect 12529 5315 12587 5321
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 13814 5312 13820 5364
rect 13872 5312 13878 5364
rect 14550 5312 14556 5364
rect 14608 5352 14614 5364
rect 14829 5355 14887 5361
rect 14829 5352 14841 5355
rect 14608 5324 14841 5352
rect 14608 5312 14614 5324
rect 14829 5321 14841 5324
rect 14875 5321 14887 5355
rect 14829 5315 14887 5321
rect 9493 5287 9551 5293
rect 9493 5253 9505 5287
rect 9539 5253 9551 5287
rect 11609 5287 11667 5293
rect 11609 5284 11621 5287
rect 11086 5256 11621 5284
rect 9493 5247 9551 5253
rect 11609 5253 11621 5256
rect 11655 5253 11667 5287
rect 11609 5247 11667 5253
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 7837 5219 7895 5225
rect 7837 5185 7849 5219
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 8021 5219 8079 5225
rect 8021 5185 8033 5219
rect 8067 5216 8079 5219
rect 8110 5216 8116 5228
rect 8067 5188 8116 5216
rect 8067 5185 8079 5188
rect 8021 5179 8079 5185
rect 7558 5108 7564 5160
rect 7616 5148 7622 5160
rect 7852 5148 7880 5179
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8481 5219 8539 5225
rect 8481 5216 8493 5219
rect 8352 5188 8493 5216
rect 8352 5176 8358 5188
rect 8481 5185 8493 5188
rect 8527 5185 8539 5219
rect 8481 5179 8539 5185
rect 8757 5219 8815 5225
rect 8757 5185 8769 5219
rect 8803 5216 8815 5219
rect 9508 5216 9536 5247
rect 8803 5188 9536 5216
rect 8803 5185 8815 5188
rect 8757 5179 8815 5185
rect 9582 5176 9588 5228
rect 9640 5176 9646 5228
rect 11698 5176 11704 5228
rect 11756 5176 11762 5228
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5216 12403 5219
rect 12434 5216 12440 5228
rect 12391 5188 12440 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12434 5176 12440 5188
rect 12492 5176 12498 5228
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 13262 5176 13268 5228
rect 13320 5216 13326 5228
rect 13357 5219 13415 5225
rect 13357 5216 13369 5219
rect 13320 5188 13369 5216
rect 13320 5176 13326 5188
rect 13357 5185 13369 5188
rect 13403 5185 13415 5219
rect 13725 5219 13783 5225
rect 13725 5216 13737 5219
rect 13357 5179 13415 5185
rect 13556 5188 13737 5216
rect 8220 5148 8248 5176
rect 7616 5120 8248 5148
rect 7616 5108 7622 5120
rect 9030 5108 9036 5160
rect 9088 5108 9094 5160
rect 9858 5108 9864 5160
rect 9916 5108 9922 5160
rect 9048 5080 9076 5108
rect 9048 5052 9352 5080
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 9033 5015 9091 5021
rect 9033 5012 9045 5015
rect 6144 4984 9045 5012
rect 6144 4972 6150 4984
rect 9033 4981 9045 4984
rect 9079 4981 9091 5015
rect 9033 4975 9091 4981
rect 9122 4972 9128 5024
rect 9180 4972 9186 5024
rect 9324 5021 9352 5052
rect 11698 5040 11704 5092
rect 11756 5080 11762 5092
rect 13556 5089 13584 5188
rect 13725 5185 13737 5188
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 14458 5176 14464 5228
rect 14516 5176 14522 5228
rect 14737 5219 14795 5225
rect 14737 5216 14749 5219
rect 14660 5188 14749 5216
rect 14660 5089 14688 5188
rect 14737 5185 14749 5188
rect 14783 5185 14795 5219
rect 14737 5179 14795 5185
rect 13541 5083 13599 5089
rect 13541 5080 13553 5083
rect 11756 5052 13553 5080
rect 11756 5040 11762 5052
rect 13541 5049 13553 5052
rect 13587 5049 13599 5083
rect 13541 5043 13599 5049
rect 14645 5083 14703 5089
rect 14645 5049 14657 5083
rect 14691 5049 14703 5083
rect 14645 5043 14703 5049
rect 9309 5015 9367 5021
rect 9309 4981 9321 5015
rect 9355 4981 9367 5015
rect 9309 4975 9367 4981
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12618 5012 12624 5024
rect 12492 4984 12624 5012
rect 12492 4972 12498 4984
rect 12618 4972 12624 4984
rect 12676 4972 12682 5024
rect 1104 4922 15456 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 15456 4922
rect 1104 4848 15456 4870
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3881 4811 3939 4817
rect 3881 4808 3893 4811
rect 3568 4780 3893 4808
rect 3568 4768 3574 4780
rect 3881 4777 3893 4780
rect 3927 4777 3939 4811
rect 3881 4771 3939 4777
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 4706 4808 4712 4820
rect 4571 4780 4712 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5442 4808 5448 4820
rect 5307 4780 5448 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5442 4768 5448 4780
rect 5500 4808 5506 4820
rect 5810 4808 5816 4820
rect 5500 4780 5816 4808
rect 5500 4768 5506 4780
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 5902 4768 5908 4820
rect 5960 4768 5966 4820
rect 7929 4811 7987 4817
rect 7929 4777 7941 4811
rect 7975 4808 7987 4811
rect 8294 4808 8300 4820
rect 7975 4780 8300 4808
rect 7975 4777 7987 4780
rect 7929 4771 7987 4777
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 9953 4811 10011 4817
rect 9953 4777 9965 4811
rect 9999 4808 10011 4811
rect 10594 4808 10600 4820
rect 9999 4780 10600 4808
rect 9999 4777 10011 4780
rect 9953 4771 10011 4777
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 4154 4700 4160 4752
rect 4212 4740 4218 4752
rect 4617 4743 4675 4749
rect 4617 4740 4629 4743
rect 4212 4712 4629 4740
rect 4212 4700 4218 4712
rect 4617 4709 4629 4712
rect 4663 4709 4675 4743
rect 4617 4703 4675 4709
rect 5077 4743 5135 4749
rect 5077 4709 5089 4743
rect 5123 4740 5135 4743
rect 5350 4740 5356 4752
rect 5123 4712 5356 4740
rect 5123 4709 5135 4712
rect 5077 4703 5135 4709
rect 5350 4700 5356 4712
rect 5408 4700 5414 4752
rect 8128 4712 9812 4740
rect 3329 4675 3387 4681
rect 3329 4641 3341 4675
rect 3375 4672 3387 4675
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 3375 4644 4353 4672
rect 3375 4641 3387 4644
rect 3329 4635 3387 4641
rect 4341 4641 4353 4644
rect 4387 4672 4399 4675
rect 4522 4672 4528 4684
rect 4387 4644 4528 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4522 4632 4528 4644
rect 4580 4672 4586 4684
rect 4798 4672 4804 4684
rect 4580 4644 4804 4672
rect 4580 4632 4586 4644
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 4985 4675 5043 4681
rect 4985 4641 4997 4675
rect 5031 4672 5043 4675
rect 5442 4672 5448 4684
rect 5031 4644 5448 4672
rect 5031 4641 5043 4644
rect 4985 4635 5043 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 3602 4564 3608 4616
rect 3660 4564 3666 4616
rect 4065 4607 4123 4613
rect 4065 4573 4077 4607
rect 4111 4573 4123 4607
rect 4065 4567 4123 4573
rect 1857 4539 1915 4545
rect 1857 4505 1869 4539
rect 1903 4505 1915 4539
rect 3513 4539 3571 4545
rect 3513 4536 3525 4539
rect 3082 4508 3525 4536
rect 1857 4499 1915 4505
rect 3513 4505 3525 4508
rect 3559 4505 3571 4539
rect 4080 4536 4108 4567
rect 4154 4564 4160 4616
rect 4212 4564 4218 4616
rect 4433 4607 4491 4613
rect 4433 4573 4445 4607
rect 4479 4604 4491 4607
rect 4706 4604 4712 4616
rect 4479 4576 4712 4604
rect 4479 4573 4491 4576
rect 4433 4567 4491 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 6178 4564 6184 4616
rect 6236 4564 6242 4616
rect 8128 4613 8156 4712
rect 9030 4672 9036 4684
rect 8404 4644 9036 4672
rect 8404 4613 8432 4644
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 9784 4672 9812 4712
rect 9858 4700 9864 4752
rect 9916 4740 9922 4752
rect 10137 4743 10195 4749
rect 10137 4740 10149 4743
rect 9916 4712 10149 4740
rect 9916 4700 9922 4712
rect 10137 4709 10149 4712
rect 10183 4709 10195 4743
rect 10137 4703 10195 4709
rect 9950 4672 9956 4684
rect 9784 4644 9956 4672
rect 8113 4607 8171 4613
rect 8113 4573 8125 4607
rect 8159 4573 8171 4607
rect 8297 4607 8355 4613
rect 8297 4604 8309 4607
rect 8113 4567 8171 4573
rect 8220 4576 8309 4604
rect 4246 4536 4252 4548
rect 4080 4508 4252 4536
rect 3513 4499 3571 4505
rect 1872 4468 1900 4499
rect 4246 4496 4252 4508
rect 4304 4496 4310 4548
rect 4798 4496 4804 4548
rect 4856 4536 4862 4548
rect 5276 4536 5304 4564
rect 5445 4539 5503 4545
rect 5445 4536 5457 4539
rect 4856 4508 5457 4536
rect 4856 4496 4862 4508
rect 5445 4505 5457 4508
rect 5491 4536 5503 4539
rect 6362 4536 6368 4548
rect 5491 4508 6368 4536
rect 5491 4505 5503 4508
rect 5445 4499 5503 4505
rect 6362 4496 6368 4508
rect 6420 4496 6426 4548
rect 6457 4539 6515 4545
rect 6457 4505 6469 4539
rect 6503 4505 6515 4539
rect 6457 4499 6515 4505
rect 2774 4468 2780 4480
rect 1872 4440 2780 4468
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 5245 4471 5303 4477
rect 5245 4437 5257 4471
rect 5291 4468 5303 4471
rect 5626 4468 5632 4480
rect 5291 4440 5632 4468
rect 5291 4437 5303 4440
rect 5245 4431 5303 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 5902 4428 5908 4480
rect 5960 4428 5966 4480
rect 6089 4471 6147 4477
rect 6089 4437 6101 4471
rect 6135 4468 6147 4471
rect 6472 4468 6500 4499
rect 7466 4496 7472 4548
rect 7524 4496 7530 4548
rect 7742 4496 7748 4548
rect 7800 4536 7806 4548
rect 8220 4536 8248 4576
rect 8297 4573 8309 4576
rect 8343 4573 8355 4607
rect 8297 4567 8355 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8481 4607 8539 4613
rect 8481 4573 8493 4607
rect 8527 4604 8539 4607
rect 8938 4604 8944 4616
rect 8527 4576 8944 4604
rect 8527 4573 8539 4576
rect 8481 4567 8539 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9048 4604 9076 4632
rect 9118 4607 9176 4613
rect 9118 4604 9130 4607
rect 9048 4576 9130 4604
rect 9118 4573 9130 4576
rect 9164 4604 9176 4607
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 9164 4576 9597 4604
rect 9164 4573 9176 4576
rect 9118 4567 9176 4573
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 9033 4539 9091 4545
rect 9033 4536 9045 4539
rect 7800 4508 9045 4536
rect 7800 4496 7806 4508
rect 9033 4505 9045 4508
rect 9079 4505 9091 4539
rect 9784 4536 9812 4644
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 13262 4632 13268 4684
rect 13320 4672 13326 4684
rect 13320 4644 14228 4672
rect 13320 4632 13326 4644
rect 12618 4564 12624 4616
rect 12676 4604 12682 4616
rect 13722 4604 13728 4616
rect 12676 4576 13728 4604
rect 12676 4564 12682 4576
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14200 4613 14228 4644
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4604 14243 4607
rect 14918 4604 14924 4616
rect 14231 4576 14924 4604
rect 14231 4573 14243 4576
rect 14185 4567 14243 4573
rect 14918 4564 14924 4576
rect 14976 4564 14982 4616
rect 9953 4539 10011 4545
rect 9953 4536 9965 4539
rect 9784 4508 9965 4536
rect 9033 4499 9091 4505
rect 9953 4505 9965 4508
rect 9999 4505 10011 4539
rect 9953 4499 10011 4505
rect 12434 4496 12440 4548
rect 12492 4496 12498 4548
rect 14458 4496 14464 4548
rect 14516 4496 14522 4548
rect 6135 4440 6500 4468
rect 6135 4437 6147 4440
rect 6089 4431 6147 4437
rect 8754 4428 8760 4480
rect 8812 4428 8818 4480
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 12805 4471 12863 4477
rect 12805 4468 12817 4471
rect 12768 4440 12817 4468
rect 12768 4428 12774 4440
rect 12805 4437 12817 4440
rect 12851 4437 12863 4471
rect 12805 4431 12863 4437
rect 1104 4378 15456 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 15456 4378
rect 1104 4304 15456 4326
rect 2774 4224 2780 4276
rect 2832 4224 2838 4276
rect 2945 4267 3003 4273
rect 2945 4233 2957 4267
rect 2991 4264 3003 4267
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 2991 4236 5365 4264
rect 2991 4233 3003 4236
rect 2945 4227 3003 4233
rect 5353 4233 5365 4236
rect 5399 4233 5411 4267
rect 5353 4227 5411 4233
rect 5442 4224 5448 4276
rect 5500 4224 5506 4276
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 5592 4236 5641 4264
rect 5592 4224 5598 4236
rect 5629 4233 5641 4236
rect 5675 4233 5687 4267
rect 5629 4227 5687 4233
rect 5902 4224 5908 4276
rect 5960 4264 5966 4276
rect 7561 4267 7619 4273
rect 7561 4264 7573 4267
rect 5960 4236 7573 4264
rect 5960 4224 5966 4236
rect 7561 4233 7573 4236
rect 7607 4233 7619 4267
rect 7561 4227 7619 4233
rect 12437 4267 12495 4273
rect 12437 4233 12449 4267
rect 12483 4264 12495 4267
rect 12729 4267 12787 4273
rect 12729 4264 12741 4267
rect 12483 4236 12741 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 12729 4233 12741 4236
rect 12775 4233 12787 4267
rect 12729 4227 12787 4233
rect 3050 4156 3056 4208
rect 3108 4196 3114 4208
rect 3145 4199 3203 4205
rect 3145 4196 3157 4199
rect 3108 4168 3157 4196
rect 3108 4156 3114 4168
rect 3145 4165 3157 4168
rect 3191 4196 3203 4199
rect 3418 4196 3424 4208
rect 3191 4168 3424 4196
rect 3191 4165 3203 4168
rect 3145 4159 3203 4165
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 4522 4196 4528 4208
rect 3528 4168 4528 4196
rect 3528 4137 3556 4168
rect 4522 4156 4528 4168
rect 4580 4196 4586 4208
rect 4617 4199 4675 4205
rect 4617 4196 4629 4199
rect 4580 4168 4629 4196
rect 4580 4156 4586 4168
rect 4617 4165 4629 4168
rect 4663 4165 4675 4199
rect 4617 4159 4675 4165
rect 4798 4156 4804 4208
rect 4856 4205 4862 4208
rect 4856 4199 4875 4205
rect 4863 4165 4875 4199
rect 5460 4196 5488 4224
rect 4856 4159 4875 4165
rect 5184 4168 5488 4196
rect 5552 4196 5580 4224
rect 6365 4199 6423 4205
rect 6365 4196 6377 4199
rect 5552 4168 6377 4196
rect 4856 4156 4862 4159
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4128 3847 4131
rect 4062 4128 4068 4140
rect 3835 4100 4068 4128
rect 3835 4097 3847 4100
rect 3789 4091 3847 4097
rect 3712 3992 3740 4091
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4246 4088 4252 4140
rect 4304 4088 4310 4140
rect 4341 4131 4399 4137
rect 4341 4097 4353 4131
rect 4387 4128 4399 4131
rect 5184 4128 5212 4168
rect 4387 4100 5212 4128
rect 5261 4131 5319 4137
rect 4387 4097 4399 4100
rect 4341 4091 4399 4097
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 5552 4128 5580 4168
rect 6365 4165 6377 4168
rect 6411 4165 6423 4199
rect 6365 4159 6423 4165
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 6549 4199 6607 4205
rect 6549 4196 6561 4199
rect 6512 4168 6561 4196
rect 6512 4156 6518 4168
rect 6549 4165 6561 4168
rect 6595 4165 6607 4199
rect 6549 4159 6607 4165
rect 8754 4156 8760 4208
rect 8812 4156 8818 4208
rect 12526 4156 12532 4208
rect 12584 4156 12590 4208
rect 14490 4168 15056 4196
rect 5491 4100 5580 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 5276 4060 5304 4091
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5684 4100 5825 4128
rect 5684 4088 5690 4100
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 5718 4060 5724 4072
rect 5000 4032 5724 4060
rect 4154 3992 4160 4004
rect 3712 3964 4160 3992
rect 4154 3952 4160 3964
rect 4212 3992 4218 4004
rect 5000 4001 5028 4032
rect 5718 4020 5724 4032
rect 5776 4020 5782 4072
rect 5828 4060 5856 4091
rect 5902 4088 5908 4140
rect 5960 4088 5966 4140
rect 6822 4088 6828 4140
rect 6880 4128 6886 4140
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 6880 4100 7205 4128
rect 6880 4088 6886 4100
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7466 4128 7472 4140
rect 7331 4100 7472 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 10413 4131 10471 4137
rect 10413 4128 10425 4131
rect 9890 4100 10425 4128
rect 10413 4097 10425 4100
rect 10459 4097 10471 4131
rect 10413 4091 10471 4097
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 11698 4128 11704 4140
rect 10551 4100 11704 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 12253 4131 12311 4137
rect 12253 4097 12265 4131
rect 12299 4128 12311 4131
rect 12342 4128 12348 4140
rect 12299 4100 12348 4128
rect 12299 4097 12311 4100
rect 12253 4091 12311 4097
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12437 4131 12495 4137
rect 12437 4097 12449 4131
rect 12483 4128 12495 4131
rect 12618 4128 12624 4140
rect 12483 4100 12624 4128
rect 12483 4097 12495 4100
rect 12437 4091 12495 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12986 4088 12992 4140
rect 13044 4088 13050 4140
rect 14550 4088 14556 4140
rect 14608 4128 14614 4140
rect 15028 4137 15056 4168
rect 14921 4131 14979 4137
rect 14921 4128 14933 4131
rect 14608 4100 14933 4128
rect 14608 4088 14614 4100
rect 14921 4097 14933 4100
rect 14967 4097 14979 4131
rect 14921 4091 14979 4097
rect 15013 4131 15071 4137
rect 15013 4097 15025 4131
rect 15059 4097 15071 4131
rect 15013 4091 15071 4097
rect 6086 4060 6092 4072
rect 5828 4032 6092 4060
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 6178 4020 6184 4072
rect 6236 4060 6242 4072
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 6236 4032 8493 4060
rect 6236 4020 6242 4032
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 8481 4023 8539 4029
rect 12912 4032 13277 4060
rect 12912 4001 12940 4032
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 13722 4020 13728 4072
rect 13780 4060 13786 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 13780 4032 14749 4060
rect 13780 4020 13786 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14737 4023 14795 4029
rect 4985 3995 5043 4001
rect 4212 3964 4660 3992
rect 4212 3952 4218 3964
rect 4632 3936 4660 3964
rect 4985 3961 4997 3995
rect 5031 3961 5043 3995
rect 4985 3955 5043 3961
rect 12897 3995 12955 4001
rect 12897 3961 12909 3995
rect 12943 3961 12955 3995
rect 12897 3955 12955 3961
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 3329 3927 3387 3933
rect 3329 3924 3341 3927
rect 3007 3896 3341 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 3329 3893 3341 3896
rect 3375 3893 3387 3927
rect 3329 3887 3387 3893
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 4801 3927 4859 3933
rect 4801 3924 4813 3927
rect 4672 3896 4813 3924
rect 4672 3884 4678 3896
rect 4801 3893 4813 3896
rect 4847 3893 4859 3927
rect 4801 3887 4859 3893
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 6733 3927 6791 3933
rect 6733 3924 6745 3927
rect 5776 3896 6745 3924
rect 5776 3884 5782 3896
rect 6733 3893 6745 3896
rect 6779 3893 6791 3927
rect 6733 3887 6791 3893
rect 8938 3884 8944 3936
rect 8996 3924 9002 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 8996 3896 10241 3924
rect 8996 3884 9002 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 12710 3884 12716 3936
rect 12768 3884 12774 3936
rect 1104 3834 15456 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 15456 3834
rect 1104 3760 15456 3782
rect 3418 3680 3424 3732
rect 3476 3720 3482 3732
rect 4430 3720 4436 3732
rect 3476 3692 4436 3720
rect 3476 3680 3482 3692
rect 4430 3680 4436 3692
rect 4488 3720 4494 3732
rect 5721 3723 5779 3729
rect 5721 3720 5733 3723
rect 4488 3692 5733 3720
rect 4488 3680 4494 3692
rect 5721 3689 5733 3692
rect 5767 3720 5779 3723
rect 5994 3720 6000 3732
rect 5767 3692 6000 3720
rect 5767 3689 5779 3692
rect 5721 3683 5779 3689
rect 5994 3680 6000 3692
rect 6052 3680 6058 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 14458 3720 14464 3732
rect 6880 3692 14464 3720
rect 6880 3680 6886 3692
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 14918 3680 14924 3732
rect 14976 3680 14982 3732
rect 4522 3652 4528 3664
rect 4172 3624 4528 3652
rect 4172 3584 4200 3624
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 5350 3612 5356 3664
rect 5408 3612 5414 3664
rect 5442 3612 5448 3664
rect 5500 3652 5506 3664
rect 6914 3652 6920 3664
rect 5500 3624 6920 3652
rect 5500 3612 5506 3624
rect 6914 3612 6920 3624
rect 6972 3612 6978 3664
rect 12526 3612 12532 3664
rect 12584 3612 12590 3664
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4080 3556 4200 3584
rect 4264 3556 4629 3584
rect 4080 3525 4108 3556
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4264 3525 4292 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4430 3476 4436 3528
rect 4488 3476 4494 3528
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3516 4767 3519
rect 5368 3516 5396 3612
rect 4755 3488 5396 3516
rect 4755 3485 4767 3488
rect 4709 3479 4767 3485
rect 4172 3448 4200 3476
rect 4724 3448 4752 3479
rect 15102 3476 15108 3528
rect 15160 3476 15166 3528
rect 4172 3420 4752 3448
rect 5718 3408 5724 3460
rect 5776 3408 5782 3460
rect 12253 3451 12311 3457
rect 12253 3417 12265 3451
rect 12299 3448 12311 3451
rect 12434 3448 12440 3460
rect 12299 3420 12440 3448
rect 12299 3417 12311 3420
rect 12253 3411 12311 3417
rect 12434 3408 12440 3420
rect 12492 3448 12498 3460
rect 13078 3448 13084 3460
rect 12492 3420 13084 3448
rect 12492 3408 12498 3420
rect 13078 3408 13084 3420
rect 13136 3408 13142 3460
rect 3789 3383 3847 3389
rect 3789 3349 3801 3383
rect 3835 3380 3847 3383
rect 4062 3380 4068 3392
rect 3835 3352 4068 3380
rect 3835 3349 3847 3352
rect 3789 3343 3847 3349
rect 4062 3340 4068 3352
rect 4120 3340 4126 3392
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 7834 3380 7840 3392
rect 5951 3352 7840 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 7834 3340 7840 3352
rect 7892 3340 7898 3392
rect 12713 3383 12771 3389
rect 12713 3349 12725 3383
rect 12759 3380 12771 3383
rect 12802 3380 12808 3392
rect 12759 3352 12808 3380
rect 12759 3349 12771 3352
rect 12713 3343 12771 3349
rect 12802 3340 12808 3352
rect 12860 3340 12866 3392
rect 1104 3290 15456 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 15456 3290
rect 1104 3216 15456 3238
rect 6178 3176 6184 3188
rect 1964 3148 6184 3176
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 1964 3049 1992 3148
rect 3234 3068 3240 3120
rect 3292 3068 3298 3120
rect 3804 3049 3832 3148
rect 6178 3136 6184 3148
rect 6236 3176 6242 3188
rect 6236 3148 8156 3176
rect 6236 3136 6242 3148
rect 4062 3068 4068 3120
rect 4120 3068 4126 3120
rect 5721 3111 5779 3117
rect 5721 3108 5733 3111
rect 5290 3080 5733 3108
rect 5721 3077 5733 3080
rect 5767 3077 5779 3111
rect 5721 3071 5779 3077
rect 7834 3068 7840 3120
rect 7892 3068 7898 3120
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1636 3012 1961 3040
rect 1636 3000 1642 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 5810 3000 5816 3052
rect 5868 3040 5874 3052
rect 5868 3012 6684 3040
rect 5868 3000 5874 3012
rect 2222 2932 2228 2984
rect 2280 2932 2286 2984
rect 4522 2932 4528 2984
rect 4580 2972 4586 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 4580 2944 5549 2972
rect 4580 2932 4586 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 6362 2932 6368 2984
rect 6420 2932 6426 2984
rect 6656 2972 6684 3012
rect 6730 3000 6736 3052
rect 6788 3000 6794 3052
rect 8128 3049 8156 3148
rect 8478 3136 8484 3188
rect 8536 3136 8542 3188
rect 12986 3136 12992 3188
rect 13044 3136 13050 3188
rect 13078 3136 13084 3188
rect 13136 3176 13142 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 13136 3148 14289 3176
rect 13136 3136 13142 3148
rect 14277 3145 14289 3148
rect 14323 3145 14335 3179
rect 14277 3139 14335 3145
rect 13004 3108 13032 3136
rect 14553 3111 14611 3117
rect 14553 3108 14565 3111
rect 12544 3080 13032 3108
rect 14030 3080 14565 3108
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 8386 3000 8392 3052
rect 8444 3000 8450 3052
rect 12544 3049 12572 3080
rect 14553 3077 14565 3080
rect 14599 3077 14611 3111
rect 14553 3071 14611 3077
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14516 3012 14657 3040
rect 14516 3000 14522 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 6822 2972 6828 2984
rect 6656 2944 6828 2972
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 12802 2932 12808 2984
rect 12860 2932 12866 2984
rect 3697 2839 3755 2845
rect 3697 2805 3709 2839
rect 3743 2836 3755 2839
rect 4614 2836 4620 2848
rect 3743 2808 4620 2836
rect 3743 2805 3755 2808
rect 3697 2799 3755 2805
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 1104 2746 15456 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 15456 2746
rect 1104 2672 15456 2694
rect 2041 2635 2099 2641
rect 2041 2601 2053 2635
rect 2087 2632 2099 2635
rect 2222 2632 2228 2644
rect 2087 2604 2228 2632
rect 2087 2601 2099 2604
rect 2041 2595 2099 2601
rect 2222 2592 2228 2604
rect 2280 2592 2286 2644
rect 3145 2635 3203 2641
rect 3145 2601 3157 2635
rect 3191 2632 3203 2635
rect 3234 2632 3240 2644
rect 3191 2604 3240 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 4706 2592 4712 2644
rect 4764 2632 4770 2644
rect 4985 2635 5043 2641
rect 4985 2632 4997 2635
rect 4764 2604 4997 2632
rect 4764 2592 4770 2604
rect 4985 2601 4997 2604
rect 5031 2601 5043 2635
rect 4985 2595 5043 2601
rect 6730 2592 6736 2644
rect 6788 2592 6794 2644
rect 6914 2592 6920 2644
rect 6972 2592 6978 2644
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8110 2632 8116 2644
rect 8067 2604 8116 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8110 2592 8116 2604
rect 8168 2592 8174 2644
rect 8386 2592 8392 2644
rect 8444 2632 8450 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 8444 2604 8493 2632
rect 8444 2592 8450 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 3050 2564 3056 2576
rect 2240 2536 3056 2564
rect 2240 2505 2268 2536
rect 3050 2524 3056 2536
rect 3108 2524 3114 2576
rect 3602 2524 3608 2576
rect 3660 2564 3666 2576
rect 5810 2564 5816 2576
rect 3660 2536 5816 2564
rect 3660 2524 3666 2536
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 7193 2567 7251 2573
rect 7193 2564 7205 2567
rect 6886 2536 7205 2564
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2465 2283 2499
rect 3789 2499 3847 2505
rect 3789 2496 3801 2499
rect 2225 2459 2283 2465
rect 2332 2468 3801 2496
rect 2332 2437 2360 2468
rect 3789 2465 3801 2468
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 4433 2499 4491 2505
rect 4433 2465 4445 2499
rect 4479 2496 4491 2499
rect 4614 2496 4620 2508
rect 4479 2468 4620 2496
rect 4479 2465 4491 2468
rect 4433 2459 4491 2465
rect 2317 2431 2375 2437
rect 2317 2397 2329 2431
rect 2363 2397 2375 2431
rect 2317 2391 2375 2397
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3602 2428 3608 2440
rect 3283 2400 3608 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3602 2388 3608 2400
rect 3660 2388 3666 2440
rect 4540 2437 4568 2468
rect 4614 2456 4620 2468
rect 4672 2456 4678 2508
rect 6886 2496 6914 2536
rect 7193 2533 7205 2536
rect 7239 2533 7251 2567
rect 7193 2527 7251 2533
rect 5092 2468 6914 2496
rect 5092 2437 5120 2468
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 5077 2431 5135 2437
rect 4571 2400 4605 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 5077 2397 5089 2431
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5810 2388 5816 2440
rect 5868 2428 5874 2440
rect 6641 2431 6699 2437
rect 6641 2428 6653 2431
rect 5868 2400 6653 2428
rect 5868 2388 5874 2400
rect 6641 2397 6653 2400
rect 6687 2397 6699 2431
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6641 2391 6699 2397
rect 6886 2400 7113 2428
rect 6454 2320 6460 2372
rect 6512 2360 6518 2372
rect 6886 2360 6914 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7190 2388 7196 2440
rect 7248 2428 7254 2440
rect 7377 2431 7435 2437
rect 7377 2428 7389 2431
rect 7248 2400 7389 2428
rect 7248 2388 7254 2400
rect 7377 2397 7389 2400
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 7837 2431 7895 2437
rect 7837 2428 7849 2431
rect 7800 2400 7849 2428
rect 7800 2388 7806 2400
rect 7837 2397 7849 2400
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 8444 2400 8677 2428
rect 8444 2388 8450 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 6512 2332 6914 2360
rect 6512 2320 6518 2332
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4709 2295 4767 2301
rect 4709 2292 4721 2295
rect 3936 2264 4721 2292
rect 3936 2252 3942 2264
rect 4709 2261 4721 2264
rect 4755 2261 4767 2295
rect 4709 2255 4767 2261
rect 1104 2202 15456 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 15456 2202
rect 1104 2128 15456 2150
<< via1 >>
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 9680 16124 9732 16176
rect 8392 16056 8444 16108
rect 9036 16056 9088 16108
rect 9772 16056 9824 16108
rect 10416 16056 10468 16108
rect 10968 16056 11020 16108
rect 11612 16056 11664 16108
rect 9956 15920 10008 15972
rect 8392 15852 8444 15904
rect 8760 15852 8812 15904
rect 9220 15852 9272 15904
rect 10048 15852 10100 15904
rect 10324 15852 10376 15904
rect 11612 15852 11664 15904
rect 11888 15895 11940 15904
rect 11888 15861 11897 15895
rect 11897 15861 11931 15895
rect 11931 15861 11940 15895
rect 11888 15852 11940 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 8576 15555 8628 15564
rect 8576 15521 8585 15555
rect 8585 15521 8619 15555
rect 8619 15521 8628 15555
rect 8576 15512 8628 15521
rect 8300 15487 8352 15496
rect 8300 15453 8309 15487
rect 8309 15453 8343 15487
rect 8343 15453 8352 15487
rect 8300 15444 8352 15453
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 8760 15444 8812 15496
rect 9312 15512 9364 15564
rect 9772 15512 9824 15564
rect 9956 15487 10008 15496
rect 9956 15453 9965 15487
rect 9965 15453 9999 15487
rect 9999 15453 10008 15487
rect 9956 15444 10008 15453
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 10324 15487 10376 15496
rect 10324 15453 10333 15487
rect 10333 15453 10367 15487
rect 10367 15453 10376 15487
rect 10324 15444 10376 15453
rect 11888 15512 11940 15564
rect 9220 15419 9272 15428
rect 9220 15385 9229 15419
rect 9229 15385 9263 15419
rect 9263 15385 9272 15419
rect 9220 15376 9272 15385
rect 11520 15487 11572 15496
rect 11520 15453 11529 15487
rect 11529 15453 11563 15487
rect 11563 15453 11572 15487
rect 11520 15444 11572 15453
rect 11612 15487 11664 15496
rect 11612 15453 11621 15487
rect 11621 15453 11655 15487
rect 11655 15453 11664 15487
rect 11612 15444 11664 15453
rect 12992 15444 13044 15496
rect 11336 15376 11388 15428
rect 8300 15308 8352 15360
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 9864 15351 9916 15360
rect 9864 15317 9873 15351
rect 9873 15317 9907 15351
rect 9907 15317 9916 15351
rect 9864 15308 9916 15317
rect 10508 15351 10560 15360
rect 10508 15317 10517 15351
rect 10517 15317 10551 15351
rect 10551 15317 10560 15351
rect 10508 15308 10560 15317
rect 11796 15351 11848 15360
rect 11796 15317 11805 15351
rect 11805 15317 11839 15351
rect 11839 15317 11848 15351
rect 11796 15308 11848 15317
rect 12716 15308 12768 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 10508 15104 10560 15156
rect 11796 15104 11848 15156
rect 12256 15104 12308 15156
rect 7288 15036 7340 15088
rect 8576 15036 8628 15088
rect 8852 15036 8904 15088
rect 8208 15011 8260 15020
rect 5264 14900 5316 14952
rect 6644 14943 6696 14952
rect 6644 14909 6653 14943
rect 6653 14909 6687 14943
rect 6687 14909 6696 14943
rect 6644 14900 6696 14909
rect 8208 14977 8217 15011
rect 8217 14977 8251 15011
rect 8251 14977 8260 15011
rect 8208 14968 8260 14977
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 9496 14968 9548 15020
rect 10048 15079 10100 15088
rect 10048 15045 10057 15079
rect 10057 15045 10091 15079
rect 10091 15045 10100 15079
rect 10048 15036 10100 15045
rect 10692 15036 10744 15088
rect 12164 15079 12216 15088
rect 12164 15045 12173 15079
rect 12173 15045 12207 15079
rect 12207 15045 12216 15079
rect 12164 15036 12216 15045
rect 10324 14968 10376 15020
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 11888 15011 11940 15020
rect 11888 14977 11897 15011
rect 11897 14977 11931 15011
rect 11931 14977 11940 15011
rect 11888 14968 11940 14977
rect 11980 14968 12032 15020
rect 14188 15104 14240 15156
rect 12716 15011 12768 15020
rect 12716 14977 12725 15011
rect 12725 14977 12759 15011
rect 12759 14977 12768 15011
rect 12716 14968 12768 14977
rect 10232 14900 10284 14952
rect 12072 14900 12124 14952
rect 9864 14832 9916 14884
rect 11796 14832 11848 14884
rect 12256 14832 12308 14884
rect 10048 14807 10100 14816
rect 10048 14773 10057 14807
rect 10057 14773 10091 14807
rect 10091 14773 10100 14807
rect 10048 14764 10100 14773
rect 10968 14764 11020 14816
rect 12348 14764 12400 14816
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 14648 14900 14700 14952
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 3976 14603 4028 14612
rect 3976 14569 3985 14603
rect 3985 14569 4019 14603
rect 4019 14569 4028 14603
rect 3976 14560 4028 14569
rect 7288 14560 7340 14612
rect 8300 14560 8352 14612
rect 11980 14560 12032 14612
rect 1676 14356 1728 14408
rect 11888 14492 11940 14544
rect 14556 14492 14608 14544
rect 10048 14424 10100 14476
rect 6000 14356 6052 14408
rect 8300 14399 8352 14408
rect 8300 14365 8309 14399
rect 8309 14365 8343 14399
rect 8343 14365 8352 14399
rect 8300 14356 8352 14365
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 3884 14288 3936 14340
rect 4712 14288 4764 14340
rect 5448 14288 5500 14340
rect 8760 14288 8812 14340
rect 9772 14288 9824 14340
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 11796 14424 11848 14476
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 2596 14220 2648 14272
rect 3792 14263 3844 14272
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 9680 14220 9732 14272
rect 11612 14220 11664 14272
rect 12256 14220 12308 14272
rect 13452 14220 13504 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 2872 13948 2924 14000
rect 5264 14016 5316 14068
rect 3792 13991 3844 14000
rect 3792 13957 3801 13991
rect 3801 13957 3835 13991
rect 3835 13957 3844 13991
rect 3792 13948 3844 13957
rect 4804 13948 4856 14000
rect 6460 13948 6512 14000
rect 6644 14016 6696 14068
rect 6920 13948 6972 14000
rect 8024 13948 8076 14000
rect 8208 13948 8260 14000
rect 10232 14016 10284 14068
rect 13268 14016 13320 14068
rect 6000 13923 6052 13932
rect 6000 13889 6009 13923
rect 6009 13889 6043 13923
rect 6043 13889 6052 13923
rect 6000 13880 6052 13889
rect 1676 13812 1728 13864
rect 2964 13855 3016 13864
rect 2964 13821 2973 13855
rect 2973 13821 3007 13855
rect 3007 13821 3016 13855
rect 2964 13812 3016 13821
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 7012 13812 7064 13864
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 8760 13923 8812 13932
rect 8760 13889 8769 13923
rect 8769 13889 8803 13923
rect 8803 13889 8812 13923
rect 8760 13880 8812 13889
rect 9864 13991 9916 14000
rect 9864 13957 9873 13991
rect 9873 13957 9907 13991
rect 9907 13957 9916 13991
rect 9864 13948 9916 13957
rect 7564 13812 7616 13864
rect 5448 13744 5500 13796
rect 4896 13676 4948 13728
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 7288 13744 7340 13796
rect 8024 13744 8076 13796
rect 9772 13744 9824 13796
rect 12164 13812 12216 13864
rect 10968 13744 11020 13796
rect 11520 13744 11572 13796
rect 14004 13812 14056 13864
rect 7104 13676 7156 13728
rect 7748 13676 7800 13728
rect 8300 13676 8352 13728
rect 8944 13719 8996 13728
rect 8944 13685 8953 13719
rect 8953 13685 8987 13719
rect 8987 13685 8996 13719
rect 8944 13676 8996 13685
rect 9956 13676 10008 13728
rect 12716 13676 12768 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2964 13472 3016 13524
rect 3976 13472 4028 13524
rect 4804 13472 4856 13524
rect 2872 13447 2924 13456
rect 2872 13413 2881 13447
rect 2881 13413 2915 13447
rect 2915 13413 2924 13447
rect 2872 13404 2924 13413
rect 3056 13404 3108 13456
rect 6000 13472 6052 13524
rect 6920 13472 6972 13524
rect 7472 13515 7524 13524
rect 7472 13481 7481 13515
rect 7481 13481 7515 13515
rect 7515 13481 7524 13515
rect 7472 13472 7524 13481
rect 9956 13472 10008 13524
rect 4344 13336 4396 13388
rect 848 13268 900 13320
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 2228 13268 2280 13277
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 1492 13132 1544 13184
rect 3056 13268 3108 13320
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 4160 13311 4212 13320
rect 4160 13277 4184 13311
rect 4184 13277 4212 13311
rect 4160 13268 4212 13277
rect 4252 13311 4304 13320
rect 4896 13336 4948 13388
rect 4252 13277 4267 13311
rect 4267 13277 4301 13311
rect 4301 13277 4304 13311
rect 4252 13268 4304 13277
rect 7012 13447 7064 13456
rect 7012 13413 7021 13447
rect 7021 13413 7055 13447
rect 7055 13413 7064 13447
rect 7012 13404 7064 13413
rect 5264 13379 5316 13388
rect 5264 13345 5273 13379
rect 5273 13345 5307 13379
rect 5307 13345 5316 13379
rect 5264 13336 5316 13345
rect 5540 13379 5592 13388
rect 5540 13345 5549 13379
rect 5549 13345 5583 13379
rect 5583 13345 5592 13379
rect 5540 13336 5592 13345
rect 7564 13404 7616 13456
rect 8208 13404 8260 13456
rect 11336 13404 11388 13456
rect 11612 13404 11664 13456
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 9772 13336 9824 13345
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 2780 13200 2832 13252
rect 6092 13200 6144 13252
rect 7748 13311 7800 13320
rect 7748 13277 7757 13311
rect 7757 13277 7791 13311
rect 7791 13277 7800 13311
rect 7748 13268 7800 13277
rect 8944 13268 8996 13320
rect 9496 13311 9548 13320
rect 9496 13277 9505 13311
rect 9505 13277 9539 13311
rect 9539 13277 9548 13311
rect 9496 13268 9548 13277
rect 11520 13311 11572 13320
rect 11520 13277 11529 13311
rect 11529 13277 11563 13311
rect 11563 13277 11572 13311
rect 11520 13268 11572 13277
rect 11888 13268 11940 13320
rect 11980 13268 12032 13320
rect 8024 13200 8076 13252
rect 3884 13132 3936 13184
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 14648 13515 14700 13524
rect 14648 13481 14657 13515
rect 14657 13481 14691 13515
rect 14691 13481 14700 13515
rect 14648 13472 14700 13481
rect 12716 13447 12768 13456
rect 12716 13413 12725 13447
rect 12725 13413 12759 13447
rect 12759 13413 12768 13447
rect 12716 13404 12768 13413
rect 12900 13268 12952 13320
rect 13268 13268 13320 13320
rect 14832 13311 14884 13320
rect 14832 13277 14841 13311
rect 14841 13277 14875 13311
rect 14875 13277 14884 13311
rect 14832 13268 14884 13277
rect 15200 13268 15252 13320
rect 12532 13175 12584 13184
rect 12532 13141 12541 13175
rect 12541 13141 12575 13175
rect 12575 13141 12584 13175
rect 12532 13132 12584 13141
rect 14924 13175 14976 13184
rect 14924 13141 14933 13175
rect 14933 13141 14967 13175
rect 14967 13141 14976 13175
rect 14924 13132 14976 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 1492 12903 1544 12912
rect 1492 12869 1501 12903
rect 1501 12869 1535 12903
rect 1535 12869 1544 12903
rect 1492 12860 1544 12869
rect 1860 12860 1912 12912
rect 2780 12860 2832 12912
rect 8208 12860 8260 12912
rect 9864 12928 9916 12980
rect 10968 12928 11020 12980
rect 11704 12928 11756 12980
rect 9956 12860 10008 12912
rect 12072 12860 12124 12912
rect 1860 12699 1912 12708
rect 1860 12665 1869 12699
rect 1869 12665 1903 12699
rect 1903 12665 1912 12699
rect 1860 12656 1912 12665
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 2872 12724 2924 12776
rect 11336 12792 11388 12844
rect 7472 12724 7524 12776
rect 9496 12767 9548 12776
rect 9496 12733 9505 12767
rect 9505 12733 9539 12767
rect 9539 12733 9548 12767
rect 9496 12724 9548 12733
rect 2688 12588 2740 12640
rect 3240 12631 3292 12640
rect 3240 12597 3249 12631
rect 3249 12597 3283 12631
rect 3283 12597 3292 12631
rect 3240 12588 3292 12597
rect 7472 12631 7524 12640
rect 7472 12597 7481 12631
rect 7481 12597 7515 12631
rect 7515 12597 7524 12631
rect 7472 12588 7524 12597
rect 7748 12631 7800 12640
rect 7748 12597 7757 12631
rect 7757 12597 7791 12631
rect 7791 12597 7800 12631
rect 7748 12588 7800 12597
rect 9772 12588 9824 12640
rect 11612 12724 11664 12776
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 13820 12860 13872 12912
rect 14188 12903 14240 12912
rect 14188 12869 14197 12903
rect 14197 12869 14231 12903
rect 14231 12869 14240 12903
rect 14188 12860 14240 12869
rect 13268 12792 13320 12844
rect 14648 12860 14700 12912
rect 14924 12860 14976 12912
rect 12256 12724 12308 12776
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 11336 12656 11388 12708
rect 13268 12656 13320 12708
rect 12716 12631 12768 12640
rect 12716 12597 12725 12631
rect 12725 12597 12759 12631
rect 12759 12597 12768 12631
rect 12716 12588 12768 12597
rect 12900 12631 12952 12640
rect 12900 12597 12909 12631
rect 12909 12597 12943 12631
rect 12943 12597 12952 12631
rect 12900 12588 12952 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 2596 12427 2648 12436
rect 2596 12393 2605 12427
rect 2605 12393 2639 12427
rect 2639 12393 2648 12427
rect 2596 12384 2648 12393
rect 4712 12384 4764 12436
rect 7472 12384 7524 12436
rect 8208 12384 8260 12436
rect 11612 12427 11664 12436
rect 11612 12393 11621 12427
rect 11621 12393 11655 12427
rect 11655 12393 11664 12427
rect 11612 12384 11664 12393
rect 13820 12384 13872 12436
rect 1768 12316 1820 12368
rect 2320 12316 2372 12368
rect 2688 12291 2740 12300
rect 2688 12257 2697 12291
rect 2697 12257 2731 12291
rect 2731 12257 2740 12291
rect 2688 12248 2740 12257
rect 3884 12291 3936 12300
rect 3884 12257 3893 12291
rect 3893 12257 3927 12291
rect 3927 12257 3936 12291
rect 3884 12248 3936 12257
rect 4620 12248 4672 12300
rect 5264 12248 5316 12300
rect 848 12180 900 12232
rect 2412 12180 2464 12232
rect 3424 12223 3476 12232
rect 3424 12189 3433 12223
rect 3433 12189 3467 12223
rect 3467 12189 3476 12223
rect 3424 12180 3476 12189
rect 1676 12155 1728 12164
rect 1676 12121 1685 12155
rect 1685 12121 1719 12155
rect 1719 12121 1728 12155
rect 1676 12112 1728 12121
rect 2044 12112 2096 12164
rect 2872 12112 2924 12164
rect 3056 12155 3108 12164
rect 3056 12121 3065 12155
rect 3065 12121 3099 12155
rect 3099 12121 3108 12155
rect 3056 12112 3108 12121
rect 4804 12180 4856 12232
rect 6184 12180 6236 12232
rect 6920 12223 6972 12232
rect 6920 12189 6929 12223
rect 6929 12189 6963 12223
rect 6963 12189 6972 12223
rect 6920 12180 6972 12189
rect 8760 12248 8812 12300
rect 9220 12248 9272 12300
rect 14556 12384 14608 12436
rect 7472 12180 7524 12232
rect 7748 12180 7800 12232
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 9404 12180 9456 12232
rect 9496 12223 9548 12232
rect 9496 12189 9505 12223
rect 9505 12189 9539 12223
rect 9539 12189 9548 12223
rect 9496 12180 9548 12189
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 14372 12223 14424 12232
rect 14372 12189 14381 12223
rect 14381 12189 14415 12223
rect 14415 12189 14424 12223
rect 14372 12180 14424 12189
rect 2780 12044 2832 12096
rect 4436 12087 4488 12096
rect 4436 12053 4445 12087
rect 4445 12053 4479 12087
rect 4479 12053 4488 12087
rect 4436 12044 4488 12053
rect 7196 12044 7248 12096
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 8944 12112 8996 12164
rect 11244 12112 11296 12164
rect 11888 12112 11940 12164
rect 11980 12155 12032 12164
rect 11980 12121 11989 12155
rect 11989 12121 12023 12155
rect 12023 12121 12032 12155
rect 11980 12112 12032 12121
rect 12440 12155 12492 12164
rect 12440 12121 12449 12155
rect 12449 12121 12483 12155
rect 12483 12121 12492 12155
rect 12440 12112 12492 12121
rect 13820 12112 13872 12164
rect 14280 12112 14332 12164
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 2872 11840 2924 11892
rect 3884 11840 3936 11892
rect 4436 11840 4488 11892
rect 1768 11815 1820 11824
rect 1768 11781 1777 11815
rect 1777 11781 1811 11815
rect 1811 11781 1820 11815
rect 1768 11772 1820 11781
rect 848 11704 900 11756
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2363 11747
rect 2363 11713 2372 11747
rect 2320 11704 2372 11713
rect 3240 11772 3292 11824
rect 2780 11747 2832 11756
rect 2780 11713 2789 11747
rect 2789 11713 2823 11747
rect 2823 11713 2832 11747
rect 2780 11704 2832 11713
rect 3056 11747 3108 11756
rect 3056 11713 3065 11747
rect 3065 11713 3099 11747
rect 3099 11713 3108 11747
rect 3056 11704 3108 11713
rect 3240 11636 3292 11688
rect 4344 11815 4396 11824
rect 4344 11781 4353 11815
rect 4353 11781 4387 11815
rect 4387 11781 4396 11815
rect 4344 11772 4396 11781
rect 4620 11772 4672 11824
rect 6184 11883 6236 11892
rect 6184 11849 6193 11883
rect 6193 11849 6227 11883
rect 6227 11849 6236 11883
rect 6184 11840 6236 11849
rect 7196 11883 7248 11892
rect 7196 11849 7205 11883
rect 7205 11849 7239 11883
rect 7239 11849 7248 11883
rect 7196 11840 7248 11849
rect 9220 11883 9272 11892
rect 9220 11849 9229 11883
rect 9229 11849 9263 11883
rect 9263 11849 9272 11883
rect 9220 11840 9272 11849
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 12072 11883 12124 11892
rect 12072 11849 12081 11883
rect 12081 11849 12115 11883
rect 12115 11849 12124 11883
rect 12072 11840 12124 11849
rect 12256 11883 12308 11892
rect 7288 11772 7340 11824
rect 9772 11815 9824 11824
rect 9772 11781 9781 11815
rect 9781 11781 9815 11815
rect 9815 11781 9824 11815
rect 9772 11772 9824 11781
rect 10508 11772 10560 11824
rect 6552 11747 6604 11756
rect 6552 11713 6561 11747
rect 6561 11713 6595 11747
rect 6595 11713 6604 11747
rect 6552 11704 6604 11713
rect 4712 11636 4764 11688
rect 2044 11611 2096 11620
rect 2044 11577 2053 11611
rect 2053 11577 2087 11611
rect 2087 11577 2096 11611
rect 2044 11568 2096 11577
rect 5816 11568 5868 11620
rect 8668 11704 8720 11756
rect 8760 11704 8812 11756
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 12256 11849 12283 11883
rect 12283 11849 12308 11883
rect 12256 11840 12308 11849
rect 12992 11840 13044 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 12532 11815 12584 11824
rect 12532 11781 12541 11815
rect 12541 11781 12575 11815
rect 12575 11781 12584 11815
rect 12532 11772 12584 11781
rect 9036 11636 9088 11688
rect 9496 11679 9548 11688
rect 9496 11645 9505 11679
rect 9505 11645 9539 11679
rect 9539 11645 9548 11679
rect 9496 11636 9548 11645
rect 11888 11636 11940 11688
rect 14004 11704 14056 11756
rect 14648 11747 14700 11756
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 12440 11568 12492 11620
rect 2320 11500 2372 11552
rect 2780 11500 2832 11552
rect 6184 11500 6236 11552
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 7196 11543 7248 11552
rect 7196 11509 7205 11543
rect 7205 11509 7239 11543
rect 7239 11509 7248 11543
rect 7196 11500 7248 11509
rect 7288 11500 7340 11552
rect 11704 11500 11756 11552
rect 12716 11543 12768 11552
rect 12716 11509 12725 11543
rect 12725 11509 12759 11543
rect 12759 11509 12768 11543
rect 12716 11500 12768 11509
rect 14372 11500 14424 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 2320 11296 2372 11348
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 3056 11228 3108 11280
rect 3240 11160 3292 11212
rect 2504 10956 2556 11008
rect 3424 11092 3476 11144
rect 4252 11296 4304 11348
rect 4896 11296 4948 11348
rect 8760 11339 8812 11348
rect 8760 11305 8769 11339
rect 8769 11305 8803 11339
rect 8803 11305 8812 11339
rect 8760 11296 8812 11305
rect 10508 11339 10560 11348
rect 10508 11305 10517 11339
rect 10517 11305 10551 11339
rect 10551 11305 10560 11339
rect 10508 11296 10560 11305
rect 4620 11228 4672 11280
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 4804 11160 4856 11212
rect 7288 11203 7340 11212
rect 7288 11169 7297 11203
rect 7297 11169 7331 11203
rect 7331 11169 7340 11203
rect 7288 11160 7340 11169
rect 14004 11296 14056 11348
rect 14924 11339 14976 11348
rect 14924 11305 14933 11339
rect 14933 11305 14967 11339
rect 14967 11305 14976 11339
rect 14924 11296 14976 11305
rect 4896 11092 4948 11144
rect 6460 11092 6512 11144
rect 7012 11135 7064 11144
rect 7012 11101 7021 11135
rect 7021 11101 7055 11135
rect 7055 11101 7064 11135
rect 7012 11092 7064 11101
rect 9312 11092 9364 11144
rect 9404 11092 9456 11144
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 11796 11092 11848 11144
rect 11980 11135 12032 11144
rect 11980 11101 11989 11135
rect 11989 11101 12023 11135
rect 12023 11101 12032 11135
rect 11980 11092 12032 11101
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12256 11092 12308 11144
rect 4804 11024 4856 11076
rect 13636 11067 13688 11076
rect 13636 11033 13645 11067
rect 13645 11033 13679 11067
rect 13679 11033 13688 11067
rect 13636 11024 13688 11033
rect 14188 11067 14240 11076
rect 14188 11033 14197 11067
rect 14197 11033 14231 11067
rect 14231 11033 14240 11067
rect 14188 11024 14240 11033
rect 15108 11135 15160 11144
rect 15108 11101 15117 11135
rect 15117 11101 15151 11135
rect 15151 11101 15160 11135
rect 15108 11092 15160 11101
rect 15200 11024 15252 11076
rect 3884 10956 3936 11008
rect 11888 10956 11940 11008
rect 12256 10956 12308 11008
rect 14280 10956 14332 11008
rect 14740 10956 14792 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 4712 10752 4764 10804
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 4068 10684 4120 10736
rect 4252 10727 4304 10736
rect 4252 10693 4261 10727
rect 4261 10693 4295 10727
rect 4295 10693 4304 10727
rect 4252 10684 4304 10693
rect 10140 10727 10192 10736
rect 10140 10693 10149 10727
rect 10149 10693 10183 10727
rect 10183 10693 10192 10727
rect 10140 10684 10192 10693
rect 12532 10752 12584 10804
rect 14188 10684 14240 10736
rect 14372 10727 14424 10736
rect 14372 10693 14381 10727
rect 14381 10693 14415 10727
rect 14415 10693 14424 10727
rect 14372 10684 14424 10693
rect 14464 10727 14516 10736
rect 14464 10693 14473 10727
rect 14473 10693 14507 10727
rect 14507 10693 14516 10727
rect 14464 10684 14516 10693
rect 848 10616 900 10668
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 2872 10616 2924 10668
rect 3240 10548 3292 10600
rect 6000 10616 6052 10668
rect 7288 10616 7340 10668
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 10508 10659 10560 10668
rect 10508 10625 10517 10659
rect 10517 10625 10551 10659
rect 10551 10625 10560 10659
rect 10508 10616 10560 10625
rect 11244 10616 11296 10668
rect 11704 10616 11756 10668
rect 12164 10659 12216 10668
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 14280 10659 14332 10668
rect 7472 10548 7524 10600
rect 9404 10548 9456 10600
rect 14280 10625 14289 10659
rect 14289 10625 14323 10659
rect 14323 10625 14332 10659
rect 14280 10616 14332 10625
rect 14648 10659 14700 10668
rect 14648 10625 14657 10659
rect 14657 10625 14691 10659
rect 14691 10625 14700 10659
rect 14648 10616 14700 10625
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 3056 10480 3108 10532
rect 3884 10523 3936 10532
rect 3884 10489 3893 10523
rect 3893 10489 3927 10523
rect 3927 10489 3936 10523
rect 3884 10480 3936 10489
rect 3148 10455 3200 10464
rect 3148 10421 3157 10455
rect 3157 10421 3191 10455
rect 3191 10421 3200 10455
rect 3148 10412 3200 10421
rect 3792 10455 3844 10464
rect 3792 10421 3801 10455
rect 3801 10421 3835 10455
rect 3835 10421 3844 10455
rect 3792 10412 3844 10421
rect 5264 10412 5316 10464
rect 6920 10412 6972 10464
rect 9312 10412 9364 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 10324 10455 10376 10464
rect 10324 10421 10333 10455
rect 10333 10421 10367 10455
rect 10367 10421 10376 10455
rect 10324 10412 10376 10421
rect 11888 10455 11940 10464
rect 11888 10421 11897 10455
rect 11897 10421 11931 10455
rect 11931 10421 11940 10455
rect 11888 10412 11940 10421
rect 14004 10412 14056 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 9956 10208 10008 10260
rect 11704 10251 11756 10260
rect 11704 10217 11713 10251
rect 11713 10217 11747 10251
rect 11747 10217 11756 10251
rect 11704 10208 11756 10217
rect 12072 10208 12124 10260
rect 2044 10140 2096 10192
rect 5632 10140 5684 10192
rect 11980 10140 12032 10192
rect 4620 10072 4672 10124
rect 5540 10072 5592 10124
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 7288 10072 7340 10124
rect 9036 10115 9088 10124
rect 9036 10081 9045 10115
rect 9045 10081 9079 10115
rect 9079 10081 9088 10115
rect 9036 10072 9088 10081
rect 9312 10115 9364 10124
rect 9312 10081 9321 10115
rect 9321 10081 9355 10115
rect 9355 10081 9364 10115
rect 9312 10072 9364 10081
rect 10508 10072 10560 10124
rect 6368 10004 6420 10056
rect 1768 9936 1820 9988
rect 1952 9911 2004 9920
rect 1952 9877 1961 9911
rect 1961 9877 1995 9911
rect 1995 9877 2004 9911
rect 1952 9868 2004 9877
rect 4620 9936 4672 9988
rect 5264 9936 5316 9988
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 6828 10004 6880 10056
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 12072 10072 12124 10124
rect 12256 10183 12308 10192
rect 12256 10149 12265 10183
rect 12265 10149 12299 10183
rect 12299 10149 12308 10183
rect 12256 10140 12308 10149
rect 13452 10251 13504 10260
rect 13452 10217 13461 10251
rect 13461 10217 13495 10251
rect 13495 10217 13504 10251
rect 13452 10208 13504 10217
rect 14648 10208 14700 10260
rect 11244 10047 11296 10056
rect 11244 10013 11253 10047
rect 11253 10013 11287 10047
rect 11287 10013 11296 10047
rect 14004 10072 14056 10124
rect 11244 10004 11296 10013
rect 9312 9936 9364 9988
rect 10324 9936 10376 9988
rect 11796 9936 11848 9988
rect 12256 9936 12308 9988
rect 7104 9868 7156 9920
rect 11060 9868 11112 9920
rect 11980 9911 12032 9920
rect 11980 9877 11989 9911
rect 11989 9877 12023 9911
rect 12023 9877 12032 9911
rect 11980 9868 12032 9877
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 14280 10047 14332 10056
rect 14280 10013 14289 10047
rect 14289 10013 14323 10047
rect 14323 10013 14332 10047
rect 14280 10004 14332 10013
rect 14188 9936 14240 9988
rect 14464 10004 14516 10056
rect 15108 10047 15160 10056
rect 15108 10013 15117 10047
rect 15117 10013 15151 10047
rect 15151 10013 15160 10047
rect 15108 10004 15160 10013
rect 13820 9911 13872 9920
rect 13820 9877 13829 9911
rect 13829 9877 13863 9911
rect 13863 9877 13872 9911
rect 13820 9868 13872 9877
rect 14924 9911 14976 9920
rect 14924 9877 14933 9911
rect 14933 9877 14967 9911
rect 14967 9877 14976 9911
rect 14924 9868 14976 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 2044 9528 2096 9580
rect 2504 9571 2556 9580
rect 2504 9537 2513 9571
rect 2513 9537 2547 9571
rect 2547 9537 2556 9571
rect 2504 9528 2556 9537
rect 3056 9571 3108 9580
rect 3056 9537 3065 9571
rect 3065 9537 3099 9571
rect 3099 9537 3108 9571
rect 3056 9528 3108 9537
rect 2320 9503 2372 9512
rect 2320 9469 2329 9503
rect 2329 9469 2363 9503
rect 2363 9469 2372 9503
rect 2320 9460 2372 9469
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 1768 9435 1820 9444
rect 1768 9401 1777 9435
rect 1777 9401 1811 9435
rect 1811 9401 1820 9435
rect 1768 9392 1820 9401
rect 4620 9664 4672 9716
rect 12532 9664 12584 9716
rect 14280 9664 14332 9716
rect 3976 9528 4028 9580
rect 4896 9528 4948 9580
rect 7288 9596 7340 9648
rect 7380 9639 7432 9648
rect 7380 9605 7389 9639
rect 7389 9605 7423 9639
rect 7423 9605 7432 9639
rect 7380 9596 7432 9605
rect 8944 9639 8996 9648
rect 8944 9605 8953 9639
rect 8953 9605 8987 9639
rect 8987 9605 8996 9639
rect 8944 9596 8996 9605
rect 9312 9639 9364 9648
rect 9312 9605 9321 9639
rect 9321 9605 9355 9639
rect 9355 9605 9364 9639
rect 9312 9596 9364 9605
rect 10140 9639 10192 9648
rect 10140 9605 10149 9639
rect 10149 9605 10183 9639
rect 10183 9605 10192 9639
rect 10140 9596 10192 9605
rect 5632 9528 5684 9580
rect 6460 9571 6512 9580
rect 6460 9537 6469 9571
rect 6469 9537 6503 9571
rect 6503 9537 6512 9571
rect 6460 9528 6512 9537
rect 9404 9571 9456 9580
rect 9404 9537 9413 9571
rect 9413 9537 9447 9571
rect 9447 9537 9456 9571
rect 9404 9528 9456 9537
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 10876 9528 10928 9580
rect 1952 9324 2004 9376
rect 4620 9392 4672 9444
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 5172 9503 5224 9512
rect 5172 9469 5181 9503
rect 5181 9469 5215 9503
rect 5215 9469 5224 9503
rect 5172 9460 5224 9469
rect 6276 9392 6328 9444
rect 2780 9324 2832 9376
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 3148 9367 3200 9376
rect 3148 9333 3157 9367
rect 3157 9333 3191 9367
rect 3191 9333 3200 9367
rect 3148 9324 3200 9333
rect 7196 9460 7248 9512
rect 11244 9528 11296 9580
rect 12256 9571 12308 9580
rect 12256 9537 12265 9571
rect 12265 9537 12299 9571
rect 12299 9537 12308 9571
rect 12256 9528 12308 9537
rect 12348 9528 12400 9580
rect 14464 9596 14516 9648
rect 13452 9528 13504 9580
rect 14648 9571 14700 9580
rect 14648 9537 14657 9571
rect 14657 9537 14691 9571
rect 14691 9537 14700 9571
rect 14648 9528 14700 9537
rect 14924 9571 14976 9580
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 11428 9460 11480 9512
rect 11888 9460 11940 9512
rect 14188 9460 14240 9512
rect 12440 9392 12492 9444
rect 11520 9324 11572 9376
rect 12072 9324 12124 9376
rect 13176 9324 13228 9376
rect 13360 9324 13412 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2504 9120 2556 9172
rect 2136 9095 2188 9104
rect 2136 9061 2145 9095
rect 2145 9061 2179 9095
rect 2179 9061 2188 9095
rect 2136 9052 2188 9061
rect 2780 9052 2832 9104
rect 2964 9163 3016 9172
rect 2964 9129 2973 9163
rect 2973 9129 3007 9163
rect 3007 9129 3016 9163
rect 2964 9120 3016 9129
rect 4620 9120 4672 9172
rect 4804 9120 4856 9172
rect 6368 9120 6420 9172
rect 3148 8984 3200 9036
rect 848 8916 900 8968
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 2688 8916 2740 8968
rect 2872 8916 2924 8968
rect 3332 8916 3384 8968
rect 5080 9052 5132 9104
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 4804 8984 4856 9036
rect 4988 8984 5040 9036
rect 5356 8984 5408 9036
rect 4896 8959 4948 8968
rect 4896 8925 4905 8959
rect 4905 8925 4939 8959
rect 4939 8925 4948 8959
rect 4896 8916 4948 8925
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5724 8959 5776 8968
rect 5724 8925 5733 8959
rect 5733 8925 5767 8959
rect 5767 8925 5776 8959
rect 5724 8916 5776 8925
rect 7012 8984 7064 9036
rect 9404 9052 9456 9104
rect 13452 9120 13504 9172
rect 14648 9120 14700 9172
rect 10508 8984 10560 9036
rect 5632 8848 5684 8900
rect 1860 8780 1912 8832
rect 2044 8780 2096 8832
rect 3976 8780 4028 8832
rect 4528 8780 4580 8832
rect 5080 8780 5132 8832
rect 5264 8780 5316 8832
rect 8484 8916 8536 8968
rect 9680 8916 9732 8968
rect 9772 8959 9824 8968
rect 9772 8925 9781 8959
rect 9781 8925 9815 8959
rect 9815 8925 9824 8959
rect 9772 8916 9824 8925
rect 11704 8984 11756 9036
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 10876 8916 10928 8968
rect 11888 8959 11940 8968
rect 11888 8925 11897 8959
rect 11897 8925 11931 8959
rect 11931 8925 11940 8959
rect 11888 8916 11940 8925
rect 15108 8984 15160 9036
rect 14188 8916 14240 8968
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 7564 8848 7616 8900
rect 6644 8780 6696 8832
rect 11428 8848 11480 8900
rect 12348 8848 12400 8900
rect 13176 8848 13228 8900
rect 14464 8891 14516 8900
rect 14464 8857 14473 8891
rect 14473 8857 14507 8891
rect 14507 8857 14516 8891
rect 14464 8848 14516 8857
rect 12164 8780 12216 8832
rect 14004 8780 14056 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2320 8576 2372 8628
rect 2688 8576 2740 8628
rect 4620 8576 4672 8628
rect 5264 8576 5316 8628
rect 5724 8576 5776 8628
rect 2136 8508 2188 8560
rect 3056 8508 3108 8560
rect 1400 8483 1452 8492
rect 1400 8449 1409 8483
rect 1409 8449 1443 8483
rect 1443 8449 1452 8483
rect 1400 8440 1452 8449
rect 1952 8440 2004 8492
rect 4528 8440 4580 8492
rect 5080 8440 5132 8492
rect 5356 8508 5408 8560
rect 6552 8576 6604 8628
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 7564 8576 7616 8628
rect 11336 8619 11388 8628
rect 11336 8585 11345 8619
rect 11345 8585 11379 8619
rect 11379 8585 11388 8619
rect 11336 8576 11388 8585
rect 11520 8576 11572 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 14648 8576 14700 8628
rect 5448 8440 5500 8492
rect 5816 8440 5868 8492
rect 2780 8372 2832 8424
rect 3332 8372 3384 8424
rect 3884 8372 3936 8424
rect 4620 8372 4672 8424
rect 5632 8415 5684 8424
rect 5632 8381 5641 8415
rect 5641 8381 5675 8415
rect 5675 8381 5684 8415
rect 5632 8372 5684 8381
rect 6644 8440 6696 8492
rect 6920 8440 6972 8492
rect 8484 8551 8536 8560
rect 8484 8517 8493 8551
rect 8493 8517 8527 8551
rect 8527 8517 8536 8551
rect 8484 8508 8536 8517
rect 10600 8508 10652 8560
rect 12164 8508 12216 8560
rect 13452 8551 13504 8560
rect 13452 8517 13461 8551
rect 13461 8517 13495 8551
rect 13495 8517 13504 8551
rect 13452 8508 13504 8517
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 7748 8483 7800 8492
rect 7748 8449 7757 8483
rect 7757 8449 7791 8483
rect 7791 8449 7800 8483
rect 7748 8440 7800 8449
rect 6460 8372 6512 8424
rect 13268 8440 13320 8492
rect 13636 8440 13688 8492
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 14280 8483 14332 8492
rect 14280 8449 14289 8483
rect 14289 8449 14323 8483
rect 14323 8449 14332 8483
rect 14280 8440 14332 8449
rect 14740 8440 14792 8492
rect 15108 8483 15160 8492
rect 15108 8449 15117 8483
rect 15117 8449 15151 8483
rect 15151 8449 15160 8483
rect 15108 8440 15160 8449
rect 1860 8347 1912 8356
rect 1860 8313 1869 8347
rect 1869 8313 1903 8347
rect 1903 8313 1912 8347
rect 1860 8304 1912 8313
rect 2872 8304 2924 8356
rect 9588 8415 9640 8424
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 1676 8236 1728 8288
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 6276 8236 6328 8288
rect 11428 8236 11480 8288
rect 11796 8236 11848 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 4712 8032 4764 8084
rect 5080 8075 5132 8084
rect 5080 8041 5089 8075
rect 5089 8041 5123 8075
rect 5123 8041 5132 8075
rect 5080 8032 5132 8041
rect 5356 8032 5408 8084
rect 5632 8032 5684 8084
rect 5908 8032 5960 8084
rect 7748 8032 7800 8084
rect 8760 8032 8812 8084
rect 3240 7964 3292 8016
rect 848 7828 900 7880
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 4804 7896 4856 7948
rect 2228 7828 2280 7837
rect 2044 7760 2096 7812
rect 2688 7760 2740 7812
rect 3700 7828 3752 7880
rect 5356 7939 5408 7948
rect 5356 7905 5365 7939
rect 5365 7905 5399 7939
rect 5399 7905 5408 7939
rect 5356 7896 5408 7905
rect 9404 7964 9456 8016
rect 9772 8032 9824 8084
rect 9956 8032 10008 8084
rect 9864 7964 9916 8016
rect 10600 8032 10652 8084
rect 11428 8032 11480 8084
rect 14280 8032 14332 8084
rect 14740 8032 14792 8084
rect 11796 7964 11848 8016
rect 7932 7828 7984 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 8852 7828 8904 7880
rect 4988 7760 5040 7812
rect 5264 7760 5316 7812
rect 9404 7803 9456 7812
rect 9404 7769 9438 7803
rect 9438 7769 9456 7803
rect 9404 7760 9456 7769
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 1860 7692 1912 7701
rect 2136 7735 2188 7744
rect 2136 7701 2145 7735
rect 2145 7701 2179 7735
rect 2179 7701 2188 7735
rect 2136 7692 2188 7701
rect 3240 7735 3292 7744
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 3516 7692 3568 7744
rect 5724 7735 5776 7744
rect 5724 7701 5733 7735
rect 5733 7701 5767 7735
rect 5767 7701 5776 7735
rect 5724 7692 5776 7701
rect 7840 7692 7892 7744
rect 9128 7692 9180 7744
rect 9772 7828 9824 7880
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 13360 7896 13412 7948
rect 9864 7692 9916 7744
rect 10876 7803 10928 7812
rect 10876 7769 10885 7803
rect 10885 7769 10919 7803
rect 10919 7769 10928 7803
rect 10876 7760 10928 7769
rect 11336 7828 11388 7880
rect 14464 7964 14516 8016
rect 14648 7896 14700 7948
rect 11796 7760 11848 7812
rect 13728 7760 13780 7812
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 15108 7871 15160 7880
rect 15108 7837 15117 7871
rect 15117 7837 15151 7871
rect 15151 7837 15160 7871
rect 15108 7828 15160 7837
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 2136 7420 2188 7472
rect 1584 7352 1636 7404
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 2872 7395 2924 7404
rect 2872 7361 2881 7395
rect 2881 7361 2915 7395
rect 2915 7361 2924 7395
rect 2872 7352 2924 7361
rect 3700 7531 3752 7540
rect 3700 7497 3709 7531
rect 3709 7497 3743 7531
rect 3743 7497 3752 7531
rect 3700 7488 3752 7497
rect 5724 7531 5776 7540
rect 5724 7497 5733 7531
rect 5733 7497 5767 7531
rect 5767 7497 5776 7531
rect 5724 7488 5776 7497
rect 3792 7463 3844 7472
rect 3792 7429 3801 7463
rect 3801 7429 3835 7463
rect 3835 7429 3844 7463
rect 3792 7420 3844 7429
rect 4804 7420 4856 7472
rect 7932 7488 7984 7540
rect 9128 7531 9180 7540
rect 9128 7497 9137 7531
rect 9137 7497 9171 7531
rect 9171 7497 9180 7531
rect 9128 7488 9180 7497
rect 7840 7463 7892 7472
rect 7840 7429 7849 7463
rect 7849 7429 7883 7463
rect 7883 7429 7892 7463
rect 7840 7420 7892 7429
rect 8392 7463 8444 7472
rect 8392 7429 8409 7463
rect 8409 7429 8444 7463
rect 8392 7420 8444 7429
rect 9956 7420 10008 7472
rect 3884 7352 3936 7404
rect 3976 7395 4028 7404
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 5356 7395 5408 7404
rect 5356 7361 5365 7395
rect 5365 7361 5399 7395
rect 5399 7361 5408 7395
rect 5356 7352 5408 7361
rect 6736 7352 6788 7404
rect 8484 7395 8536 7404
rect 8484 7361 8493 7395
rect 8493 7361 8527 7395
rect 8527 7361 8536 7395
rect 8484 7352 8536 7361
rect 2228 7284 2280 7336
rect 1676 7216 1728 7268
rect 3240 7216 3292 7268
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 3332 7191 3384 7200
rect 3332 7157 3341 7191
rect 3341 7157 3375 7191
rect 3375 7157 3384 7191
rect 3332 7148 3384 7157
rect 8208 7327 8260 7336
rect 8208 7293 8217 7327
rect 8217 7293 8251 7327
rect 8251 7293 8260 7327
rect 8208 7284 8260 7293
rect 9128 7352 9180 7404
rect 8852 7284 8904 7336
rect 9588 7352 9640 7404
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 9772 7216 9824 7268
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 9588 7148 9640 7200
rect 11796 7148 11848 7200
rect 13176 7148 13228 7200
rect 13728 7148 13780 7200
rect 14372 7148 14424 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 3976 6944 4028 6996
rect 5356 6944 5408 6996
rect 6000 6944 6052 6996
rect 8300 6944 8352 6996
rect 8484 6944 8536 6996
rect 11704 6987 11756 6996
rect 11704 6953 11713 6987
rect 11713 6953 11747 6987
rect 11747 6953 11756 6987
rect 11704 6944 11756 6953
rect 11980 6944 12032 6996
rect 12164 6944 12216 6996
rect 1584 6876 1636 6928
rect 1952 6808 2004 6860
rect 2780 6808 2832 6860
rect 5448 6808 5500 6860
rect 6736 6808 6788 6860
rect 8208 6876 8260 6928
rect 10876 6876 10928 6928
rect 4252 6740 4304 6792
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 7564 6740 7616 6792
rect 8760 6808 8812 6860
rect 9312 6851 9364 6860
rect 9312 6817 9321 6851
rect 9321 6817 9355 6851
rect 9355 6817 9364 6851
rect 9312 6808 9364 6817
rect 9128 6740 9180 6792
rect 12716 6740 12768 6792
rect 12992 6783 13044 6792
rect 12992 6749 13001 6783
rect 13001 6749 13035 6783
rect 13035 6749 13044 6783
rect 12992 6740 13044 6749
rect 6092 6672 6144 6724
rect 6920 6672 6972 6724
rect 8944 6672 8996 6724
rect 12440 6672 12492 6724
rect 13176 6783 13228 6792
rect 13176 6749 13185 6783
rect 13185 6749 13219 6783
rect 13219 6749 13228 6783
rect 13176 6740 13228 6749
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 13728 6740 13780 6792
rect 14372 6783 14424 6792
rect 14372 6749 14381 6783
rect 14381 6749 14415 6783
rect 14415 6749 14424 6783
rect 14372 6740 14424 6749
rect 5724 6647 5776 6656
rect 5724 6613 5751 6647
rect 5751 6613 5776 6647
rect 5724 6604 5776 6613
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 9680 6604 9732 6613
rect 12992 6604 13044 6656
rect 13452 6604 13504 6656
rect 13636 6647 13688 6656
rect 13636 6613 13645 6647
rect 13645 6613 13679 6647
rect 13679 6613 13688 6647
rect 13636 6604 13688 6613
rect 13728 6647 13780 6656
rect 13728 6613 13737 6647
rect 13737 6613 13771 6647
rect 13771 6613 13780 6647
rect 13728 6604 13780 6613
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14556 6672 14608 6724
rect 15108 6783 15160 6792
rect 15108 6749 15117 6783
rect 15117 6749 15151 6783
rect 15151 6749 15160 6783
rect 15108 6740 15160 6749
rect 14924 6647 14976 6656
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2688 6400 2740 6452
rect 4620 6400 4672 6452
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 9312 6400 9364 6452
rect 848 6264 900 6316
rect 4068 6332 4120 6384
rect 5632 6375 5684 6384
rect 5632 6341 5641 6375
rect 5641 6341 5675 6375
rect 5675 6341 5684 6375
rect 5632 6332 5684 6341
rect 9036 6332 9088 6384
rect 14188 6400 14240 6452
rect 3516 6264 3568 6316
rect 4896 6307 4948 6316
rect 4896 6273 4905 6307
rect 4905 6273 4939 6307
rect 4939 6273 4948 6307
rect 4896 6264 4948 6273
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5356 6264 5408 6316
rect 6736 6264 6788 6316
rect 8208 6264 8260 6316
rect 9128 6307 9180 6316
rect 9128 6273 9137 6307
rect 9137 6273 9171 6307
rect 9171 6273 9180 6307
rect 9128 6264 9180 6273
rect 12992 6332 13044 6384
rect 11612 6264 11664 6316
rect 11796 6264 11848 6316
rect 2872 6171 2924 6180
rect 2872 6137 2881 6171
rect 2881 6137 2915 6171
rect 2915 6137 2924 6171
rect 2872 6128 2924 6137
rect 4252 6171 4304 6180
rect 4252 6137 4261 6171
rect 4261 6137 4295 6171
rect 4295 6137 4304 6171
rect 4252 6128 4304 6137
rect 4620 6128 4672 6180
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 5264 6060 5316 6112
rect 5908 6060 5960 6112
rect 6092 6060 6144 6112
rect 6828 6060 6880 6112
rect 8576 6196 8628 6248
rect 8760 6239 8812 6248
rect 8760 6205 8769 6239
rect 8769 6205 8803 6239
rect 8803 6205 8812 6239
rect 8760 6196 8812 6205
rect 8852 6239 8904 6248
rect 8852 6205 8861 6239
rect 8861 6205 8895 6239
rect 8895 6205 8904 6239
rect 8852 6196 8904 6205
rect 11060 6239 11112 6248
rect 11060 6205 11069 6239
rect 11069 6205 11103 6239
rect 11103 6205 11112 6239
rect 11060 6196 11112 6205
rect 12440 6307 12492 6316
rect 12440 6273 12449 6307
rect 12449 6273 12483 6307
rect 12483 6273 12492 6307
rect 12440 6264 12492 6273
rect 14096 6332 14148 6384
rect 12624 6196 12676 6248
rect 13820 6307 13872 6316
rect 13820 6273 13829 6307
rect 13829 6273 13863 6307
rect 13863 6273 13872 6307
rect 13820 6264 13872 6273
rect 14372 6332 14424 6384
rect 14280 6307 14332 6316
rect 14280 6273 14289 6307
rect 14289 6273 14323 6307
rect 14323 6273 14332 6307
rect 14280 6264 14332 6273
rect 14556 6307 14608 6316
rect 14556 6273 14565 6307
rect 14565 6273 14599 6307
rect 14599 6273 14608 6307
rect 14556 6264 14608 6273
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 15200 6196 15252 6248
rect 9496 6103 9548 6112
rect 9496 6069 9505 6103
rect 9505 6069 9539 6103
rect 9539 6069 9548 6103
rect 9496 6060 9548 6069
rect 9956 6060 10008 6112
rect 12164 6128 12216 6180
rect 14740 6128 14792 6180
rect 11980 6060 12032 6112
rect 13728 6060 13780 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3884 5856 3936 5908
rect 4620 5856 4672 5908
rect 5632 5856 5684 5908
rect 8392 5856 8444 5908
rect 3056 5788 3108 5840
rect 4712 5720 4764 5772
rect 5724 5788 5776 5840
rect 5908 5788 5960 5840
rect 9680 5788 9732 5840
rect 6000 5720 6052 5772
rect 4804 5652 4856 5704
rect 4988 5652 5040 5704
rect 5448 5652 5500 5704
rect 2872 5584 2924 5636
rect 6092 5652 6144 5704
rect 6184 5652 6236 5704
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 8944 5652 8996 5704
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 11060 5856 11112 5908
rect 11888 5899 11940 5908
rect 11888 5865 11897 5899
rect 11897 5865 11931 5899
rect 11931 5865 11940 5899
rect 11888 5856 11940 5865
rect 12072 5856 12124 5908
rect 12532 5856 12584 5908
rect 13820 5856 13872 5908
rect 14556 5856 14608 5908
rect 13728 5788 13780 5840
rect 11704 5720 11756 5772
rect 12992 5720 13044 5772
rect 8484 5584 8536 5636
rect 8852 5584 8904 5636
rect 4620 5516 4672 5568
rect 4896 5516 4948 5568
rect 8760 5516 8812 5568
rect 8944 5516 8996 5568
rect 9496 5584 9548 5636
rect 10508 5584 10560 5636
rect 12072 5652 12124 5704
rect 13728 5652 13780 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 14372 5695 14424 5704
rect 14372 5661 14381 5695
rect 14381 5661 14415 5695
rect 14415 5661 14424 5695
rect 14372 5652 14424 5661
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 11980 5584 12032 5636
rect 10600 5559 10652 5568
rect 10600 5525 10609 5559
rect 10609 5525 10643 5559
rect 10643 5525 10652 5559
rect 10600 5516 10652 5525
rect 13820 5584 13872 5636
rect 12624 5516 12676 5568
rect 13360 5516 13412 5568
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 6736 5312 6788 5364
rect 8300 5312 8352 5364
rect 9036 5312 9088 5364
rect 9128 5312 9180 5364
rect 8576 5244 8628 5296
rect 8944 5244 8996 5296
rect 9772 5312 9824 5364
rect 10508 5312 10560 5364
rect 11888 5312 11940 5364
rect 13728 5312 13780 5364
rect 13820 5355 13872 5364
rect 13820 5321 13829 5355
rect 13829 5321 13863 5355
rect 13863 5321 13872 5355
rect 13820 5312 13872 5321
rect 14556 5312 14608 5364
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 7564 5108 7616 5160
rect 8116 5176 8168 5228
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 12440 5176 12492 5228
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 13268 5176 13320 5228
rect 9036 5108 9088 5160
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 6092 4972 6144 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 11704 5040 11756 5092
rect 14464 5219 14516 5228
rect 14464 5185 14473 5219
rect 14473 5185 14507 5219
rect 14507 5185 14516 5219
rect 14464 5176 14516 5185
rect 12440 4972 12492 5024
rect 12624 4972 12676 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 3516 4768 3568 4820
rect 4712 4768 4764 4820
rect 5448 4768 5500 4820
rect 5816 4768 5868 4820
rect 5908 4811 5960 4820
rect 5908 4777 5917 4811
rect 5917 4777 5951 4811
rect 5951 4777 5960 4811
rect 5908 4768 5960 4777
rect 8300 4768 8352 4820
rect 10600 4768 10652 4820
rect 4160 4700 4212 4752
rect 5356 4700 5408 4752
rect 4528 4632 4580 4684
rect 4804 4632 4856 4684
rect 5448 4632 5500 4684
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 3608 4607 3660 4616
rect 3608 4573 3617 4607
rect 3617 4573 3651 4607
rect 3651 4573 3660 4607
rect 3608 4564 3660 4573
rect 4160 4607 4212 4616
rect 4160 4573 4169 4607
rect 4169 4573 4203 4607
rect 4203 4573 4212 4607
rect 4160 4564 4212 4573
rect 4712 4564 4764 4616
rect 5264 4564 5316 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 6184 4607 6236 4616
rect 6184 4573 6193 4607
rect 6193 4573 6227 4607
rect 6227 4573 6236 4607
rect 6184 4564 6236 4573
rect 9036 4632 9088 4684
rect 9864 4700 9916 4752
rect 4252 4496 4304 4548
rect 4804 4496 4856 4548
rect 6368 4496 6420 4548
rect 2780 4428 2832 4480
rect 5632 4428 5684 4480
rect 5908 4471 5960 4480
rect 5908 4437 5917 4471
rect 5917 4437 5951 4471
rect 5951 4437 5960 4471
rect 5908 4428 5960 4437
rect 7472 4496 7524 4548
rect 7748 4496 7800 4548
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 9956 4632 10008 4684
rect 13268 4632 13320 4684
rect 12624 4607 12676 4616
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 13728 4564 13780 4616
rect 14924 4564 14976 4616
rect 12440 4539 12492 4548
rect 12440 4505 12449 4539
rect 12449 4505 12483 4539
rect 12483 4505 12492 4539
rect 12440 4496 12492 4505
rect 14464 4539 14516 4548
rect 14464 4505 14473 4539
rect 14473 4505 14507 4539
rect 14507 4505 14516 4539
rect 14464 4496 14516 4505
rect 8760 4471 8812 4480
rect 8760 4437 8769 4471
rect 8769 4437 8803 4471
rect 8803 4437 8812 4471
rect 8760 4428 8812 4437
rect 12716 4428 12768 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 2780 4267 2832 4276
rect 2780 4233 2789 4267
rect 2789 4233 2823 4267
rect 2823 4233 2832 4267
rect 2780 4224 2832 4233
rect 5448 4224 5500 4276
rect 5540 4224 5592 4276
rect 5908 4224 5960 4276
rect 3056 4156 3108 4208
rect 3424 4156 3476 4208
rect 4528 4156 4580 4208
rect 4804 4199 4856 4208
rect 4804 4165 4829 4199
rect 4829 4165 4856 4199
rect 4804 4156 4856 4165
rect 4068 4088 4120 4140
rect 4252 4131 4304 4140
rect 4252 4097 4261 4131
rect 4261 4097 4295 4131
rect 4295 4097 4304 4131
rect 4252 4088 4304 4097
rect 6460 4156 6512 4208
rect 8760 4199 8812 4208
rect 8760 4165 8769 4199
rect 8769 4165 8803 4199
rect 8803 4165 8812 4199
rect 8760 4156 8812 4165
rect 12532 4199 12584 4208
rect 12532 4165 12541 4199
rect 12541 4165 12575 4199
rect 12575 4165 12584 4199
rect 12532 4156 12584 4165
rect 5632 4088 5684 4140
rect 4160 3952 4212 4004
rect 5724 4020 5776 4072
rect 5908 4131 5960 4140
rect 5908 4097 5917 4131
rect 5917 4097 5951 4131
rect 5951 4097 5960 4131
rect 5908 4088 5960 4097
rect 6828 4088 6880 4140
rect 7472 4088 7524 4140
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 11704 4088 11756 4140
rect 12348 4088 12400 4140
rect 12624 4088 12676 4140
rect 12992 4131 13044 4140
rect 12992 4097 13001 4131
rect 13001 4097 13035 4131
rect 13035 4097 13044 4131
rect 12992 4088 13044 4097
rect 14556 4088 14608 4140
rect 6092 4020 6144 4072
rect 6184 4020 6236 4072
rect 13728 4020 13780 4072
rect 4620 3884 4672 3936
rect 5724 3884 5776 3936
rect 8944 3884 8996 3936
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3424 3680 3476 3732
rect 4436 3680 4488 3732
rect 6000 3680 6052 3732
rect 6828 3680 6880 3732
rect 14464 3680 14516 3732
rect 14924 3723 14976 3732
rect 14924 3689 14933 3723
rect 14933 3689 14967 3723
rect 14967 3689 14976 3723
rect 14924 3680 14976 3689
rect 4528 3612 4580 3664
rect 5356 3655 5408 3664
rect 5356 3621 5365 3655
rect 5365 3621 5399 3655
rect 5399 3621 5408 3655
rect 5356 3612 5408 3621
rect 5448 3612 5500 3664
rect 6920 3612 6972 3664
rect 12532 3655 12584 3664
rect 12532 3621 12541 3655
rect 12541 3621 12575 3655
rect 12575 3621 12584 3655
rect 12532 3612 12584 3621
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4436 3519 4488 3528
rect 4436 3485 4445 3519
rect 4445 3485 4479 3519
rect 4479 3485 4488 3519
rect 4436 3476 4488 3485
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 5724 3451 5776 3460
rect 5724 3417 5733 3451
rect 5733 3417 5767 3451
rect 5767 3417 5776 3451
rect 5724 3408 5776 3417
rect 12440 3408 12492 3460
rect 13084 3408 13136 3460
rect 4068 3340 4120 3392
rect 7840 3340 7892 3392
rect 12808 3340 12860 3392
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1584 3000 1636 3052
rect 3240 3068 3292 3120
rect 6184 3136 6236 3188
rect 4068 3111 4120 3120
rect 4068 3077 4077 3111
rect 4077 3077 4111 3111
rect 4111 3077 4120 3111
rect 4068 3068 4120 3077
rect 7840 3111 7892 3120
rect 7840 3077 7849 3111
rect 7849 3077 7883 3111
rect 7883 3077 7892 3111
rect 7840 3068 7892 3077
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 2228 2975 2280 2984
rect 2228 2941 2237 2975
rect 2237 2941 2271 2975
rect 2271 2941 2280 2975
rect 2228 2932 2280 2941
rect 4528 2932 4580 2984
rect 6368 2975 6420 2984
rect 6368 2941 6377 2975
rect 6377 2941 6411 2975
rect 6411 2941 6420 2975
rect 6368 2932 6420 2941
rect 6736 3000 6788 3052
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 12992 3136 13044 3188
rect 13084 3136 13136 3188
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 14464 3000 14516 3052
rect 6828 2932 6880 2984
rect 12808 2975 12860 2984
rect 12808 2941 12817 2975
rect 12817 2941 12851 2975
rect 12851 2941 12860 2975
rect 12808 2932 12860 2941
rect 4620 2796 4672 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 2228 2592 2280 2644
rect 3240 2592 3292 2644
rect 4712 2592 4764 2644
rect 6736 2635 6788 2644
rect 6736 2601 6745 2635
rect 6745 2601 6779 2635
rect 6779 2601 6788 2635
rect 6736 2592 6788 2601
rect 6920 2635 6972 2644
rect 6920 2601 6929 2635
rect 6929 2601 6963 2635
rect 6963 2601 6972 2635
rect 6920 2592 6972 2601
rect 8116 2592 8168 2644
rect 8392 2592 8444 2644
rect 3056 2524 3108 2576
rect 3608 2524 3660 2576
rect 5816 2524 5868 2576
rect 3608 2388 3660 2440
rect 4620 2456 4672 2508
rect 5816 2388 5868 2440
rect 6460 2320 6512 2372
rect 7196 2388 7248 2440
rect 7748 2388 7800 2440
rect 8392 2388 8444 2440
rect 3884 2252 3936 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 8390 17950 8446 18750
rect 9034 17950 9090 18750
rect 9678 17950 9734 18750
rect 10322 17950 10378 18750
rect 10966 17950 11022 18750
rect 11610 17950 11666 18750
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 8404 16114 8432 17950
rect 9048 16114 9076 17950
rect 9692 16182 9720 17950
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 10336 16130 10364 17950
rect 10336 16114 10456 16130
rect 10980 16114 11008 17950
rect 11624 16114 11652 17950
rect 8392 16108 8444 16114
rect 8392 16050 8444 16056
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9772 16108 9824 16114
rect 10336 16108 10468 16114
rect 10336 16102 10416 16108
rect 9772 16050 9824 16056
rect 10416 16050 10468 16056
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 8404 15502 8432 15846
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8300 15496 8352 15502
rect 8300 15438 8352 15444
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 8312 15366 8340 15438
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7378 15056 7434 15065
rect 5264 14952 5316 14958
rect 5264 14894 5316 14900
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 13870 1716 14350
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 3792 14272 3844 14278
rect 3792 14214 3844 14220
rect 1676 13864 1728 13870
rect 1676 13806 1728 13812
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 13161 888 13262
rect 1492 13184 1544 13190
rect 846 13152 902 13161
rect 1492 13126 1544 13132
rect 846 13087 902 13096
rect 1504 12918 1532 13126
rect 1492 12912 1544 12918
rect 1492 12854 1544 12860
rect 848 12232 900 12238
rect 846 12200 848 12209
rect 900 12200 902 12209
rect 1688 12170 1716 13806
rect 2608 13326 2636 14214
rect 3804 14006 3832 14214
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 2884 13462 2912 13942
rect 2964 13864 3016 13870
rect 2964 13806 3016 13812
rect 2976 13530 3004 13806
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 3056 13456 3108 13462
rect 3056 13398 3108 13404
rect 3068 13326 3096 13398
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 1860 12912 1912 12918
rect 1860 12854 1912 12860
rect 1872 12714 1900 12854
rect 1860 12708 1912 12714
rect 1860 12650 1912 12656
rect 1768 12368 1820 12374
rect 1768 12310 1820 12316
rect 846 12135 902 12144
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1780 11830 1808 12310
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 1768 11824 1820 11830
rect 846 11792 902 11801
rect 1768 11766 1820 11772
rect 846 11727 848 11736
rect 900 11727 902 11736
rect 848 11698 900 11704
rect 2056 11626 2084 12106
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 2240 11257 2268 13262
rect 2780 13252 2832 13258
rect 2780 13194 2832 13200
rect 2792 12918 2820 13194
rect 3896 13190 3924 14282
rect 3988 13530 4016 14554
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3988 13394 4384 13410
rect 3988 13388 4396 13394
rect 3988 13382 4344 13388
rect 3988 13326 4016 13382
rect 4344 13330 4396 13336
rect 3976 13320 4028 13326
rect 4160 13320 4212 13326
rect 3976 13262 4028 13268
rect 4080 13280 4160 13308
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 2608 12442 2636 12718
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2596 12436 2648 12442
rect 2596 12378 2648 12384
rect 2320 12368 2372 12374
rect 2320 12310 2372 12316
rect 2332 11762 2360 12310
rect 2700 12306 2728 12582
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2320 11552 2372 11558
rect 2424 11540 2452 12174
rect 2884 12170 2912 12718
rect 3240 12640 3292 12646
rect 3240 12582 3292 12588
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 2780 12096 2832 12102
rect 2780 12038 2832 12044
rect 2792 11762 2820 12038
rect 2884 11898 2912 12106
rect 2872 11892 2924 11898
rect 2872 11834 2924 11840
rect 3068 11762 3096 12106
rect 3252 11830 3280 12582
rect 3884 12300 3936 12306
rect 4080 12288 4108 13280
rect 4252 13320 4304 13326
rect 4212 13280 4252 13308
rect 4160 13262 4212 13268
rect 4252 13262 4304 13268
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4724 12442 4752 14282
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5276 14074 5304 14894
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4816 13530 4844 13942
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4908 13394 4936 13670
rect 5276 13394 5304 14010
rect 5460 13802 5488 14282
rect 6012 13938 6040 14350
rect 6656 14074 6684 14894
rect 7300 14618 7328 15030
rect 7378 14991 7434 15000
rect 8208 15020 8260 15026
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6460 14000 6512 14006
rect 6460 13942 6512 13948
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5552 13394 5580 13670
rect 6012 13530 6040 13874
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 5276 12306 5304 13330
rect 3936 12260 4108 12288
rect 4620 12300 4672 12306
rect 3884 12242 3936 12248
rect 4620 12242 4672 12248
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3240 11824 3292 11830
rect 3240 11766 3292 11772
rect 2780 11756 2832 11762
rect 3056 11756 3108 11762
rect 2832 11716 2912 11744
rect 2780 11698 2832 11704
rect 2372 11512 2452 11540
rect 2780 11552 2832 11558
rect 2320 11494 2372 11500
rect 2780 11494 2832 11500
rect 2332 11354 2360 11494
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2226 11248 2282 11257
rect 2226 11183 2282 11192
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 2504 11008 2556 11014
rect 1398 10976 1454 10985
rect 2504 10950 2556 10956
rect 1398 10911 1454 10920
rect 2516 10674 2544 10950
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 860 10441 888 10610
rect 846 10432 902 10441
rect 846 10367 902 10376
rect 2044 10192 2096 10198
rect 2044 10134 2096 10140
rect 1768 9988 1820 9994
rect 1768 9930 1820 9936
rect 1780 9450 1808 9930
rect 1952 9920 2004 9926
rect 1952 9862 2004 9868
rect 1768 9444 1820 9450
rect 1768 9386 1820 9392
rect 1964 9382 1992 9862
rect 2056 9586 2084 10134
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2240 9625 2268 9998
rect 2226 9616 2282 9625
rect 2044 9580 2096 9586
rect 2226 9551 2282 9560
rect 2504 9580 2556 9586
rect 2044 9522 2096 9528
rect 2504 9522 2556 9528
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 846 9072 902 9081
rect 846 9007 902 9016
rect 860 8974 888 9007
rect 848 8968 900 8974
rect 848 8910 900 8916
rect 2056 8838 2084 9522
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 1860 8832 1912 8838
rect 1860 8774 1912 8780
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1400 8492 1452 8498
rect 1400 8434 1452 8440
rect 1412 8265 1440 8434
rect 1872 8362 1900 8774
rect 2148 8566 2176 9046
rect 2332 8974 2360 9454
rect 2516 9178 2544 9522
rect 2792 9518 2820 11494
rect 2884 10674 2912 11716
rect 3056 11698 3108 11704
rect 3068 11286 3096 11698
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3056 11280 3108 11286
rect 3108 11228 3188 11234
rect 3056 11222 3188 11228
rect 3068 11206 3188 11222
rect 3252 11218 3280 11630
rect 2872 10668 2924 10674
rect 2872 10610 2924 10616
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 3068 9586 3096 10474
rect 3160 10470 3188 11206
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 10606 3280 11154
rect 3436 11150 3464 12174
rect 3896 11898 3924 12242
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11898 4476 12038
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 4436 11892 4488 11898
rect 4436 11834 4488 11840
rect 4632 11830 4660 12242
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4344 11824 4396 11830
rect 4344 11766 4396 11772
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 4356 11540 4384 11766
rect 4080 11512 4384 11540
rect 4080 11336 4108 11512
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4252 11348 4304 11354
rect 4080 11308 4252 11336
rect 4252 11290 4304 11296
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3884 11008 3936 11014
rect 3884 10950 3936 10956
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3148 10464 3200 10470
rect 3148 10406 3200 10412
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2780 9376 2832 9382
rect 2964 9376 3016 9382
rect 2832 9324 2912 9330
rect 2780 9318 2912 9324
rect 2964 9318 3016 9324
rect 2792 9302 2912 9318
rect 2504 9172 2556 9178
rect 2504 9114 2556 9120
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2688 8968 2740 8974
rect 2688 8910 2740 8916
rect 2332 8634 2360 8910
rect 2700 8634 2728 8910
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2688 8628 2740 8634
rect 2688 8570 2740 8576
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1676 8288 1728 8294
rect 1398 8256 1454 8265
rect 1676 8230 1728 8236
rect 1398 8191 1454 8200
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 1584 7744 1636 7750
rect 846 7712 902 7721
rect 1584 7686 1636 7692
rect 846 7647 902 7656
rect 1596 7410 1624 7686
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1596 6934 1624 7346
rect 1688 7274 1716 8230
rect 1964 7886 1992 8434
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1872 7410 1900 7686
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1584 6928 1636 6934
rect 1584 6870 1636 6876
rect 1964 6866 1992 7822
rect 2044 7812 2096 7818
rect 2044 7754 2096 7760
rect 2056 7546 2084 7754
rect 2136 7744 2188 7750
rect 2136 7686 2188 7692
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2148 7478 2176 7686
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2240 7342 2268 7822
rect 2700 7818 2728 8570
rect 2792 8430 2820 9046
rect 2884 8974 2912 9302
rect 2976 9178 3004 9318
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 3068 8566 3096 9522
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 9042 3188 9318
rect 3148 9036 3200 9042
rect 3148 8978 3200 8984
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2688 7812 2740 7818
rect 2688 7754 2740 7760
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2700 6458 2728 7346
rect 2792 7206 2820 8366
rect 2872 8356 2924 8362
rect 2872 8298 2924 8304
rect 2884 7410 2912 8298
rect 3252 8022 3280 10542
rect 3896 10538 3924 10950
rect 4264 10742 4292 11290
rect 4632 11286 4660 11766
rect 4712 11688 4764 11694
rect 4712 11630 4764 11636
rect 4620 11280 4672 11286
rect 4342 11248 4398 11257
rect 4620 11222 4672 11228
rect 4342 11183 4398 11192
rect 4356 11150 4384 11183
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4068 10736 4120 10742
rect 4068 10678 4120 10684
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 3884 10532 3936 10538
rect 3884 10474 3936 10480
rect 3792 10464 3844 10470
rect 3792 10406 3844 10412
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3344 8430 3372 8910
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 2872 7404 2924 7410
rect 2872 7346 2924 7352
rect 3252 7274 3280 7686
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3344 7206 3372 8366
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 2792 6866 2820 7142
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 846 6352 902 6361
rect 3528 6322 3556 7686
rect 3712 7546 3740 7822
rect 3700 7540 3752 7546
rect 3700 7482 3752 7488
rect 3804 7478 3832 10406
rect 3976 9580 4028 9586
rect 3976 9522 4028 9528
rect 3988 8838 4016 9522
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3884 8424 3936 8430
rect 3884 8366 3936 8372
rect 3792 7472 3844 7478
rect 3792 7414 3844 7420
rect 3896 7410 3924 8366
rect 4080 7410 4108 10678
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10130 4660 11222
rect 4724 11098 4752 11630
rect 4816 11218 4844 12174
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4908 11150 4936 11290
rect 4896 11144 4948 11150
rect 4724 11082 4844 11098
rect 4896 11086 4948 11092
rect 4724 11076 4856 11082
rect 4724 11070 4804 11076
rect 4804 11018 4856 11024
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4632 9722 4660 9930
rect 4620 9716 4672 9722
rect 4620 9658 4672 9664
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4632 9178 4660 9386
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8498 4568 8774
rect 4632 8634 4660 9114
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 3516 6316 3568 6322
rect 848 6258 900 6264
rect 3516 6258 3568 6264
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2884 5642 2912 6122
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5846 3096 6054
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 3528 4826 3556 6258
rect 3896 5914 3924 7346
rect 3988 7002 4016 7346
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4080 6390 4108 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4264 6186 4292 6734
rect 4632 6458 4660 8366
rect 4724 8090 4752 10746
rect 4816 9178 4844 11018
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5276 9994 5304 10406
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5264 9988 5316 9994
rect 5264 9930 5316 9936
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4816 7954 4844 8978
rect 4908 8974 4936 9522
rect 4988 9512 5040 9518
rect 5172 9512 5224 9518
rect 4988 9454 5040 9460
rect 5092 9472 5172 9500
rect 5000 9042 5028 9454
rect 5092 9110 5120 9472
rect 5172 9454 5224 9460
rect 5080 9104 5132 9110
rect 5080 9046 5132 9052
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 4896 8968 4948 8974
rect 4896 8910 4948 8916
rect 5092 8838 5120 9046
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 8774
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5368 8566 5396 8978
rect 5552 8974 5580 10066
rect 5644 9586 5672 10134
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5644 8906 5672 9522
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5736 8634 5764 8910
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4816 7478 4844 7890
rect 5000 7818 5028 8230
rect 5092 8090 5120 8434
rect 5368 8090 5396 8502
rect 5828 8498 5856 11562
rect 6012 10674 6040 13466
rect 6104 13258 6132 13806
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 6184 12232 6236 12238
rect 6184 12174 6236 12180
rect 6196 11898 6224 12174
rect 6184 11892 6236 11898
rect 6184 11834 6236 11840
rect 6196 11558 6224 11834
rect 6472 11558 6500 13942
rect 6932 13530 6960 13942
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 6932 12238 6960 13466
rect 7024 13462 7052 13806
rect 7288 13796 7340 13802
rect 7288 13738 7340 13744
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6552 11756 6604 11762
rect 6552 11698 6604 11704
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 11257 6500 11494
rect 6458 11248 6514 11257
rect 6380 11206 6458 11234
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6380 10062 6408 11206
rect 6458 11183 6514 11192
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 10810 6500 11086
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6564 10146 6592 11698
rect 7116 11540 7144 13670
rect 7300 13326 7328 13738
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7208 11898 7236 12038
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7300 11830 7328 12038
rect 7288 11824 7340 11830
rect 7288 11766 7340 11772
rect 7196 11552 7248 11558
rect 7116 11512 7196 11540
rect 7196 11494 7248 11500
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6472 10118 6592 10146
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6472 9586 6500 10118
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6828 10056 6880 10062
rect 6932 10010 6960 10406
rect 7024 10062 7052 11086
rect 6880 10004 6960 10010
rect 6828 9998 6960 10004
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6460 9580 6512 9586
rect 6460 9522 6512 9528
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5356 8084 5408 8090
rect 5356 8026 5408 8032
rect 5368 7954 5396 8026
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 4988 7812 5040 7818
rect 4988 7754 5040 7760
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 5276 6798 5304 7754
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5368 7002 5396 7346
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 5368 6322 5396 6938
rect 5460 6866 5488 8434
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5644 8090 5672 8366
rect 6288 8294 6316 9386
rect 6368 9172 6420 9178
rect 6472 9160 6500 9522
rect 6420 9132 6500 9160
rect 6368 9114 6420 9120
rect 6472 8430 6500 9132
rect 6564 8634 6592 9998
rect 6840 9982 6960 9998
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6656 8498 6684 8774
rect 6932 8498 6960 9982
rect 7024 9042 7052 9998
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7012 9036 7064 9042
rect 7012 8978 7064 8984
rect 7116 8634 7144 9862
rect 7208 9518 7236 11494
rect 7300 11218 7328 11494
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 10130 7328 10610
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 9654 7328 10066
rect 7392 9654 7420 14991
rect 8208 14962 8260 14968
rect 8220 14006 8248 14962
rect 8312 14618 8340 15302
rect 8588 15094 8616 15506
rect 8772 15502 8800 15846
rect 8760 15496 8812 15502
rect 8760 15438 8812 15444
rect 8772 15178 8800 15438
rect 9232 15434 9260 15846
rect 9784 15570 9812 16050
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9312 15564 9364 15570
rect 9312 15506 9364 15512
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9220 15428 9272 15434
rect 9220 15370 9272 15376
rect 8772 15150 8892 15178
rect 8864 15094 8892 15150
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 9324 15026 9352 15506
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9508 15026 9536 15302
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8024 14000 8076 14006
rect 8024 13942 8076 13948
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7484 13530 7512 13874
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7484 12782 7512 13466
rect 7576 13462 7604 13806
rect 8036 13802 8064 13942
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7760 13326 7788 13670
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7760 12646 7788 13262
rect 8036 13258 8064 13738
rect 8220 13462 8248 13942
rect 8312 13734 8340 14350
rect 9784 14346 9812 15506
rect 9968 15502 9996 15914
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9876 14890 9904 15302
rect 10060 15094 10088 15846
rect 10336 15502 10364 15846
rect 11624 15502 11652 15846
rect 11900 15570 11928 15846
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11612 15496 11664 15502
rect 11612 15438 11664 15444
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10244 14958 10272 15438
rect 10336 15026 10364 15438
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 10508 15360 10560 15366
rect 10508 15302 10560 15308
rect 10520 15162 10548 15302
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10692 15088 10744 15094
rect 10692 15030 10744 15036
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 14482 10088 14758
rect 10048 14476 10100 14482
rect 10048 14418 10100 14424
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 8772 13938 8800 14282
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8300 13728 8352 13734
rect 8300 13670 8352 13676
rect 8208 13456 8260 13462
rect 8208 13398 8260 13404
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7748 12640 7800 12646
rect 7748 12582 7800 12588
rect 7484 12442 7512 12582
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7760 12238 7788 12582
rect 8036 12238 8064 13194
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8220 12442 8248 12854
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7748 12232 7800 12238
rect 7748 12174 7800 12180
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7484 10606 7512 12174
rect 8680 11762 8708 13126
rect 8772 12306 8800 13874
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8956 13326 8984 13670
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9508 12782 9536 13262
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 8760 12300 8812 12306
rect 8760 12242 8812 12248
rect 9220 12300 9272 12306
rect 9220 12242 9272 12248
rect 8944 12164 8996 12170
rect 8944 12106 8996 12112
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8772 11354 8800 11698
rect 8760 11348 8812 11354
rect 8760 11290 8812 11296
rect 7472 10600 7524 10606
rect 7472 10542 7524 10548
rect 8956 9654 8984 12106
rect 9232 11898 9260 12242
rect 9508 12238 9536 12718
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 9048 10130 9076 11630
rect 9416 11150 9444 12174
rect 9508 11694 9536 12174
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9324 10996 9352 11086
rect 9324 10968 9444 10996
rect 9416 10606 9444 10968
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9324 10130 9352 10406
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9324 9654 9352 9930
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7576 8634 7604 8842
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 8496 8566 8524 8910
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 7748 8492 7800 8498
rect 7748 8434 7800 8440
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7546 5764 7686
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 4252 6180 4304 6186
rect 4252 6122 4304 6128
rect 4620 6180 4672 6186
rect 4620 6122 4672 6128
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5914 4660 6122
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4712 5772 4764 5778
rect 4712 5714 4764 5720
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 4160 4752 4212 4758
rect 4160 4694 4212 4700
rect 4172 4622 4200 4694
rect 4528 4684 4580 4690
rect 4528 4626 4580 4632
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 4160 4616 4212 4622
rect 4160 4558 4212 4564
rect 1596 3058 1624 4558
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4282 2820 4422
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2228 2984 2280 2990
rect 2228 2926 2280 2932
rect 2240 2650 2268 2926
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 3068 2582 3096 4150
rect 3436 3738 3464 4150
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3252 2650 3280 3062
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3620 2582 3648 4558
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4080 3652 4108 4082
rect 4172 4010 4200 4558
rect 4252 4548 4304 4554
rect 4252 4490 4304 4496
rect 4264 4146 4292 4490
rect 4540 4214 4568 4626
rect 4632 4604 4660 5510
rect 4724 4826 4752 5714
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4816 4690 4844 5646
rect 4908 5574 4936 6258
rect 5000 5710 5028 6258
rect 5264 6112 5316 6118
rect 5264 6054 5316 6060
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 5276 4622 5304 6054
rect 5460 5710 5488 6802
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5644 5914 5672 6326
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5736 5846 5764 6598
rect 5920 6118 5948 8026
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5846 5948 6054
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5908 5840 5960 5846
rect 5908 5782 5960 5788
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5460 4826 5488 5646
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5356 4752 5408 4758
rect 5356 4694 5408 4700
rect 4712 4616 4764 4622
rect 4632 4576 4712 4604
rect 4712 4558 4764 4564
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4080 3624 4200 3652
rect 4172 3534 4200 3624
rect 4448 3534 4476 3674
rect 4528 3664 4580 3670
rect 4632 3652 4660 3878
rect 4580 3624 4660 3652
rect 4528 3606 4580 3612
rect 4540 3534 4568 3606
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4080 3126 4108 3334
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4540 2990 4568 3470
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 3608 2576 3660 2582
rect 3608 2518 3660 2524
rect 3620 2446 3648 2518
rect 4632 2514 4660 2790
rect 4724 2650 4752 4558
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4816 4214 4844 4490
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 5368 3670 5396 4694
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5460 4282 5488 4626
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5552 4282 5580 4558
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5460 3670 5488 4218
rect 5644 4146 5672 4422
rect 5632 4140 5684 4146
rect 5632 4082 5684 4088
rect 5736 4078 5764 5782
rect 5920 4826 5948 5782
rect 6012 5778 6040 6938
rect 6748 6866 6776 7346
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 7576 6798 7604 8434
rect 7760 8090 7788 8434
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8772 7886 8800 8026
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7852 7478 7880 7686
rect 7944 7546 7972 7822
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7840 7472 7892 7478
rect 8392 7472 8444 7478
rect 7840 7414 7892 7420
rect 8312 7420 8392 7426
rect 8312 7414 8444 7420
rect 8312 7398 8432 7414
rect 8496 7410 8524 7822
rect 8484 7404 8536 7410
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 8220 6934 8248 7278
rect 8312 7002 8340 7398
rect 8484 7346 8536 7352
rect 8496 7002 8524 7346
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8208 6928 8260 6934
rect 8208 6870 8260 6876
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6104 6118 6132 6666
rect 6736 6316 6788 6322
rect 6736 6258 6788 6264
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6000 5772 6052 5778
rect 6000 5714 6052 5720
rect 6012 5012 6040 5714
rect 6104 5710 6132 6054
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6092 5024 6144 5030
rect 6012 4984 6092 5012
rect 6092 4966 6144 4972
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5828 4128 5856 4762
rect 5920 4570 5948 4762
rect 5920 4542 6040 4570
rect 5908 4480 5960 4486
rect 5908 4422 5960 4428
rect 5920 4282 5948 4422
rect 5908 4276 5960 4282
rect 5908 4218 5960 4224
rect 5908 4140 5960 4146
rect 5828 4100 5908 4128
rect 5908 4082 5960 4088
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5736 3466 5764 3878
rect 6012 3738 6040 4542
rect 6104 4078 6132 4966
rect 6196 4622 6224 5646
rect 6748 5370 6776 6258
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6840 5710 6868 6054
rect 6828 5704 6880 5710
rect 6828 5646 6880 5652
rect 6932 5556 6960 6666
rect 8220 6458 8248 6870
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 6840 5528 6960 5556
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6840 5234 6868 5528
rect 8220 5234 8248 6258
rect 8312 5370 8340 6938
rect 8772 6866 8800 7822
rect 8864 7342 8892 7822
rect 8852 7336 8904 7342
rect 8852 7278 8904 7284
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8956 6730 8984 9590
rect 9416 9586 9444 10542
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9416 9110 9444 9522
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9692 8974 9720 14214
rect 10244 14074 10272 14894
rect 10704 14414 10732 15030
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14414 11008 14758
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9772 13796 9824 13802
rect 9772 13738 9824 13744
rect 9784 13394 9812 13738
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9876 12986 9904 13942
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 9956 13728 10008 13734
rect 9956 13670 10008 13676
rect 9968 13530 9996 13670
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9968 12918 9996 13466
rect 10980 12986 11008 13738
rect 11348 13462 11376 15370
rect 11532 14498 11560 15438
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 12716 15360 12768 15366
rect 12716 15302 12768 15308
rect 11808 15178 11836 15302
rect 11716 15162 11836 15178
rect 11716 15156 11848 15162
rect 11716 15150 11796 15156
rect 11532 14470 11652 14498
rect 11624 14278 11652 14470
rect 11716 14414 11744 15150
rect 11796 15098 11848 15104
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12164 15088 12216 15094
rect 12084 15036 12164 15042
rect 12084 15030 12216 15036
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12084 15014 12204 15030
rect 11808 14890 11836 14962
rect 11796 14884 11848 14890
rect 11796 14826 11848 14832
rect 11808 14482 11836 14826
rect 11900 14550 11928 14962
rect 11992 14618 12020 14962
rect 12084 14958 12112 15014
rect 12072 14952 12124 14958
rect 12072 14894 12124 14900
rect 12268 14890 12296 15098
rect 12728 15026 12756 15302
rect 13004 15026 13032 15438
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11796 14476 11848 14482
rect 11796 14418 11848 14424
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 12256 14272 12308 14278
rect 12360 14260 12388 14758
rect 12308 14232 12388 14260
rect 12256 14214 12308 14220
rect 11520 13796 11572 13802
rect 11520 13738 11572 13744
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 11348 12850 11376 13398
rect 11532 13326 11560 13738
rect 11624 13462 11652 14214
rect 13280 14074 13308 14962
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11348 12714 11376 12786
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11336 12708 11388 12714
rect 11336 12650 11388 12656
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9784 11830 9812 12582
rect 11624 12442 11652 12718
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11256 11898 11284 12106
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 10508 11824 10560 11830
rect 10508 11766 10560 11772
rect 10520 11354 10548 11766
rect 11612 11756 11664 11762
rect 11716 11744 11744 12922
rect 11900 12850 11928 13262
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11900 12170 11928 12786
rect 11992 12170 12020 13262
rect 12072 12912 12124 12918
rect 12072 12854 12124 12860
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11664 11716 11744 11744
rect 11612 11698 11664 11704
rect 11716 11558 11744 11716
rect 11900 11694 11928 12106
rect 11992 11898 12020 12106
rect 12084 11898 12112 12854
rect 12176 12238 12204 13806
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12728 13462 12756 13670
rect 12716 13456 12768 13462
rect 12716 13398 12768 13404
rect 13280 13326 13308 14010
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10266 9996 10406
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 10152 9654 10180 10678
rect 10428 10674 10456 11086
rect 11716 10674 11744 11494
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 9994 10364 10406
rect 10520 10130 10548 10610
rect 10508 10124 10560 10130
rect 10508 10066 10560 10072
rect 11256 10062 11284 10610
rect 11716 10266 11744 10610
rect 11704 10260 11756 10266
rect 11704 10202 11756 10208
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9704 11100 9862
rect 10980 9676 11100 9704
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10876 9580 10928 9586
rect 10980 9568 11008 9676
rect 11256 9586 11284 9998
rect 11808 9994 11836 11086
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11900 10470 11928 10950
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11992 10198 12020 11086
rect 12084 10266 12112 11086
rect 12176 10674 12204 12174
rect 12268 11898 12296 12718
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12452 11626 12480 12106
rect 12544 11830 12572 13126
rect 12912 12646 12940 13262
rect 13280 12850 13308 13262
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13280 12714 13308 12786
rect 13268 12708 13320 12714
rect 13268 12650 13320 12656
rect 12716 12640 12768 12646
rect 12716 12582 12768 12588
rect 12900 12640 12952 12646
rect 12900 12582 12952 12588
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12268 11014 12296 11086
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12072 10260 12124 10266
rect 12072 10202 12124 10208
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11992 9926 12020 10134
rect 12084 10130 12112 10202
rect 12268 10198 12296 10950
rect 12544 10810 12572 11766
rect 12728 11558 12756 12582
rect 12912 12434 12940 12582
rect 12912 12406 13032 12434
rect 13004 11898 13032 12406
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12072 10124 12124 10130
rect 12072 10066 12124 10072
rect 12084 9926 12112 10066
rect 12256 9988 12308 9994
rect 12256 9930 12308 9936
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 12268 9586 12296 9930
rect 12544 9722 12572 10746
rect 13464 10266 13492 14214
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13832 12442 13860 12854
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13832 11898 13860 12106
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 14016 11762 14044 13806
rect 14200 12918 14228 15098
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14556 14544 14608 14550
rect 14556 14486 14608 14492
rect 14188 12912 14240 12918
rect 14188 12854 14240 12860
rect 14200 12238 14228 12854
rect 14568 12442 14596 14486
rect 14660 13530 14688 14894
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14660 13410 14688 13466
rect 14660 13382 14780 13410
rect 14648 12912 14700 12918
rect 14648 12854 14700 12860
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14016 11354 14044 11698
rect 14004 11348 14056 11354
rect 14004 11290 14056 11296
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 14188 11076 14240 11082
rect 14188 11018 14240 11024
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 10928 9540 11008 9568
rect 11244 9580 11296 9586
rect 10876 9522 10928 9528
rect 11244 9522 11296 9528
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12348 9580 12400 9586
rect 12348 9522 12400 9528
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 10520 9042 10548 9522
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10888 8974 10916 9522
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 9680 8968 9732 8974
rect 9680 8910 9732 8916
rect 9772 8968 9824 8974
rect 9772 8910 9824 8916
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9404 8016 9456 8022
rect 9404 7958 9456 7964
rect 9416 7818 9444 7958
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7546 9168 7686
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9140 7410 9168 7482
rect 9600 7410 9628 8366
rect 9784 8090 9812 8910
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10612 8090 10640 8502
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 9600 7206 9628 7346
rect 9784 7274 9812 7822
rect 9876 7750 9904 7958
rect 9968 7886 9996 8026
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 9864 7744 9916 7750
rect 9864 7686 9916 7692
rect 9968 7478 9996 7822
rect 10888 7818 10916 8910
rect 11440 8906 11468 9454
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11428 8900 11480 8906
rect 11428 8842 11480 8848
rect 11336 8628 11388 8634
rect 11440 8616 11468 8842
rect 11532 8634 11560 9318
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11388 8588 11468 8616
rect 11520 8628 11572 8634
rect 11336 8570 11388 8576
rect 11520 8570 11572 8576
rect 11348 7886 11376 8570
rect 11428 8288 11480 8294
rect 11428 8230 11480 8236
rect 11440 8090 11468 8230
rect 11428 8084 11480 8090
rect 11428 8026 11480 8032
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 9956 7472 10008 7478
rect 9956 7414 10008 7420
rect 9772 7268 9824 7274
rect 9772 7210 9824 7216
rect 9588 7200 9640 7206
rect 9588 7142 9640 7148
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 5914 8432 6598
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6196 4078 6224 4558
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6380 4196 6408 4490
rect 6460 4208 6512 4214
rect 6380 4168 6460 4196
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6000 3732 6052 3738
rect 6000 3674 6052 3680
rect 5724 3460 5776 3466
rect 5724 3402 5776 3408
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 6196 3194 6224 4014
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5828 2582 5856 2994
rect 6380 2990 6408 4168
rect 6460 4150 6512 4156
rect 6840 4146 6868 5170
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7472 4548 7524 4554
rect 7472 4490 7524 4496
rect 7484 4146 7512 4490
rect 7576 4146 7604 5102
rect 7748 4548 7800 4554
rect 7748 4490 7800 4496
rect 7760 4146 7788 4490
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 6840 3738 6868 4082
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6748 2650 6776 2994
rect 6840 2990 6868 3674
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6932 2650 6960 3606
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7852 3126 7880 3334
rect 7840 3120 7892 3126
rect 7840 3062 7892 3068
rect 8128 2650 8156 5170
rect 8312 4826 8340 5170
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8496 3194 8524 5578
rect 8588 5302 8616 6190
rect 8772 5574 8800 6190
rect 8864 5642 8892 6190
rect 8956 5710 8984 6666
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5302 8984 5510
rect 9048 5370 9076 6326
rect 9140 6322 9168 6734
rect 9324 6458 9352 6802
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9140 5370 9168 6258
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5642 9536 6054
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 8576 5296 8628 5302
rect 8576 5238 8628 5244
rect 8944 5296 8996 5302
rect 8944 5238 8996 5244
rect 8956 4622 8984 5238
rect 9048 5166 9076 5306
rect 9600 5234 9628 7142
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 5846 9720 6598
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9784 5370 9812 7210
rect 10888 6934 10916 7754
rect 11716 7410 11744 8978
rect 11900 8974 11928 9454
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9178 12112 9318
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 12360 8906 12388 9522
rect 12440 9444 12492 9450
rect 12440 9386 12492 9392
rect 12452 9042 12480 9386
rect 13176 9376 13228 9382
rect 13176 9318 13228 9324
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 13188 8906 13216 9318
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 13176 8900 13228 8906
rect 13176 8842 13228 8848
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 8566 12204 8774
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11808 8022 11836 8230
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11716 7002 11744 7346
rect 11808 7206 11836 7754
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11704 6996 11756 7002
rect 11704 6938 11756 6944
rect 10876 6928 10928 6934
rect 10876 6870 10928 6876
rect 11612 6316 11664 6322
rect 11716 6304 11744 6938
rect 11808 6322 11836 7142
rect 11992 7002 12020 7278
rect 12176 7002 12204 8502
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 11664 6276 11744 6304
rect 11612 6258 11664 6264
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9968 5914 9996 6054
rect 11072 5914 11100 6190
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9128 5024 9180 5030
rect 9048 4984 9128 5012
rect 9048 4690 9076 4984
rect 9128 4966 9180 4972
rect 9876 4758 9904 5102
rect 9864 4752 9916 4758
rect 9864 4694 9916 4700
rect 9968 4690 9996 5850
rect 11716 5778 11744 6276
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 10508 5636 10560 5642
rect 10508 5578 10560 5584
rect 10520 5370 10548 5578
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10612 4826 10640 5510
rect 11704 5228 11756 5234
rect 11808 5216 11836 6258
rect 12176 6186 12204 6938
rect 13188 6798 13216 7142
rect 12716 6792 12768 6798
rect 12636 6740 12716 6746
rect 12636 6734 12768 6740
rect 12992 6792 13044 6798
rect 12992 6734 13044 6740
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 12440 6724 12492 6730
rect 12440 6666 12492 6672
rect 12636 6718 12756 6734
rect 12452 6322 12480 6666
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 11980 6112 12032 6118
rect 11980 6054 12032 6060
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11900 5370 11928 5850
rect 11992 5642 12020 6054
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 12084 5710 12112 5850
rect 12072 5704 12124 5710
rect 12072 5646 12124 5652
rect 11980 5636 12032 5642
rect 11980 5578 12032 5584
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 12452 5234 12480 6258
rect 12636 6254 12664 6718
rect 13004 6662 13032 6734
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13004 6390 13032 6598
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12624 6248 12676 6254
rect 12624 6190 12676 6196
rect 12532 5908 12584 5914
rect 12532 5850 12584 5856
rect 11756 5188 11836 5216
rect 12440 5228 12492 5234
rect 11704 5170 11756 5176
rect 12440 5170 12492 5176
rect 11716 5098 11744 5170
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8760 4480 8812 4486
rect 8760 4422 8812 4428
rect 8772 4214 8800 4422
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8956 3942 8984 4558
rect 11716 4146 11744 5034
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12452 4554 12480 4966
rect 12440 4548 12492 4554
rect 12440 4490 12492 4496
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 12348 4140 12400 4146
rect 12452 4128 12480 4490
rect 12544 4214 12572 5850
rect 12636 5574 12664 6190
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12636 5234 12664 5510
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12636 5030 12664 5170
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12532 4208 12584 4214
rect 12532 4150 12584 4156
rect 12400 4100 12480 4128
rect 12348 4082 12400 4088
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 12452 3466 12480 4100
rect 12544 3670 12572 4150
rect 12636 4146 12664 4558
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12728 3942 12756 4422
rect 13004 4146 13032 5714
rect 13280 5234 13308 8434
rect 13372 7954 13400 9318
rect 13464 9178 13492 9522
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13464 8566 13492 9114
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13648 8498 13676 11018
rect 14200 10742 14228 11018
rect 14292 11014 14320 12106
rect 14384 11558 14412 12174
rect 14568 11898 14596 12174
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14660 11762 14688 12854
rect 14752 12850 14780 13382
rect 14832 13320 14884 13326
rect 14832 13262 14884 13268
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 14844 13025 14872 13262
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14830 13016 14886 13025
rect 14830 12951 14886 12960
rect 14936 12918 14964 13126
rect 14924 12912 14976 12918
rect 14924 12854 14976 12860
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 15212 12345 15240 13262
rect 15198 12336 15254 12345
rect 15198 12271 15254 12280
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14292 10674 14320 10950
rect 14384 10742 14412 11494
rect 14936 11354 14964 11698
rect 15106 11656 15162 11665
rect 15106 11591 15162 11600
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15120 11150 15148 11591
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 14740 11008 14792 11014
rect 15212 10985 15240 11018
rect 14740 10950 14792 10956
rect 15198 10976 15254 10985
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14016 10130 14044 10406
rect 14004 10124 14056 10130
rect 14004 10066 14056 10072
rect 14476 10062 14504 10678
rect 14752 10674 14780 10950
rect 15198 10911 15254 10920
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14660 10266 14688 10610
rect 15106 10296 15162 10305
rect 14648 10260 14700 10266
rect 15106 10231 15162 10240
rect 14648 10202 14700 10208
rect 15120 10062 15148 10231
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 8634 13860 9862
rect 14200 9518 14228 9930
rect 14292 9722 14320 9998
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14280 9716 14332 9722
rect 14332 9676 14412 9704
rect 14280 9658 14332 9664
rect 14188 9512 14240 9518
rect 14188 9454 14240 9460
rect 14200 8974 14228 9454
rect 14384 8974 14412 9676
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14476 8906 14504 9590
rect 14936 9586 14964 9862
rect 15106 9616 15162 9625
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14924 9580 14976 9586
rect 15106 9551 15162 9560
rect 14924 9522 14976 9528
rect 14660 9178 14688 9522
rect 14648 9172 14700 9178
rect 14648 9114 14700 9120
rect 15120 9042 15148 9551
rect 15108 9036 15160 9042
rect 15108 8978 15160 8984
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 15106 8936 15162 8945
rect 14464 8900 14516 8906
rect 14464 8842 14516 8848
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 14016 8498 14044 8774
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14280 8492 14332 8498
rect 14280 8434 14332 8440
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13740 7206 13768 7754
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 6798 13768 7142
rect 13544 6792 13596 6798
rect 13372 6740 13544 6746
rect 13372 6734 13596 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13372 6718 13584 6734
rect 13372 5574 13400 6718
rect 13452 6656 13504 6662
rect 13636 6656 13688 6662
rect 13504 6604 13636 6610
rect 13452 6598 13688 6604
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 13464 6582 13676 6598
rect 13648 5658 13676 6582
rect 13740 6118 13768 6598
rect 14108 6390 14136 6598
rect 14200 6458 14228 8434
rect 14292 8090 14320 8434
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14476 8022 14504 8842
rect 14660 8634 14688 8910
rect 15106 8871 15162 8880
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14660 7954 14688 8570
rect 15120 8498 15148 8871
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14752 8090 14780 8434
rect 15106 8256 15162 8265
rect 15106 8191 15162 8200
rect 14740 8084 14792 8090
rect 14740 8026 14792 8032
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 15120 7886 15148 8191
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 14476 7698 14504 7822
rect 14384 7670 14504 7698
rect 14384 7206 14412 7670
rect 14462 7576 14518 7585
rect 14462 7511 14518 7520
rect 14476 7410 14504 7511
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6798 14412 7142
rect 15106 6896 15162 6905
rect 15106 6831 15162 6840
rect 15120 6798 15148 6831
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 14556 6724 14608 6730
rect 14556 6666 14608 6672
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 13820 6316 13872 6322
rect 13820 6258 13872 6264
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 13728 6112 13780 6118
rect 13728 6054 13780 6060
rect 13740 5846 13768 6054
rect 13832 5914 13860 6258
rect 13820 5908 13872 5914
rect 13820 5850 13872 5856
rect 13728 5840 13780 5846
rect 13728 5782 13780 5788
rect 14292 5710 14320 6258
rect 14384 5710 14412 6326
rect 14568 6322 14596 6666
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14936 6322 14964 6598
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14924 6316 14976 6322
rect 14924 6258 14976 6264
rect 14568 5914 14596 6258
rect 15200 6248 15252 6254
rect 15198 6216 15200 6225
rect 15252 6216 15254 6225
rect 14740 6180 14792 6186
rect 15198 6151 15254 6160
rect 14740 6122 14792 6128
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 14752 5710 14780 6122
rect 13728 5704 13780 5710
rect 13648 5652 13728 5658
rect 13648 5646 13780 5652
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14372 5704 14424 5710
rect 14372 5646 14424 5652
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 13648 5630 13768 5646
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13740 5370 13768 5630
rect 13820 5636 13872 5642
rect 13820 5578 13872 5584
rect 13832 5370 13860 5578
rect 14462 5536 14518 5545
rect 14462 5471 14518 5480
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13820 5364 13872 5370
rect 13820 5306 13872 5312
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13280 4690 13308 5170
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 13740 4622 13768 5306
rect 14476 5234 14504 5471
rect 14568 5370 14596 5646
rect 14556 5364 14608 5370
rect 14556 5306 14608 5312
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 12992 4140 13044 4146
rect 12992 4082 13044 4088
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8404 2650 8432 2994
rect 12820 2990 12848 3334
rect 13004 3194 13032 4082
rect 13740 4078 13768 4558
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14476 4128 14504 4490
rect 14556 4140 14608 4146
rect 14476 4100 14556 4128
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 14476 3738 14504 4100
rect 14556 4082 14608 4088
rect 14936 3738 14964 4558
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 13084 3460 13136 3466
rect 13084 3402 13136 3408
rect 13096 3194 13124 3402
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 14476 3058 14504 3674
rect 15108 3528 15160 3534
rect 15106 3496 15108 3505
rect 15160 3496 15162 3505
rect 15106 3431 15162 3440
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 12808 2984 12860 2990
rect 12808 2926 12860 2932
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 8116 2644 8168 2650
rect 8116 2586 8168 2592
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 5828 2446 5856 2518
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 800 3924 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 6472 800 6500 2314
rect 7208 1306 7236 2382
rect 7116 1278 7236 1306
rect 7116 800 7144 1278
rect 7760 800 7788 2382
rect 8404 800 8432 2382
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
<< via2 >>
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 846 13096 902 13152
rect 846 12180 848 12200
rect 848 12180 900 12200
rect 900 12180 902 12200
rect 846 12144 902 12180
rect 846 11756 902 11792
rect 846 11736 848 11756
rect 848 11736 900 11756
rect 900 11736 902 11756
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 7378 15000 7434 15056
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 2226 11192 2282 11248
rect 1398 10920 1454 10976
rect 846 10376 902 10432
rect 2226 9560 2282 9616
rect 846 9016 902 9072
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1398 8200 1454 8256
rect 846 7656 902 7712
rect 4342 11192 4398 11248
rect 846 6316 902 6352
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 6458 11192 6514 11248
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 14830 12960 14886 13016
rect 15198 12280 15254 12336
rect 15106 11600 15162 11656
rect 15198 10920 15254 10976
rect 15106 10240 15162 10296
rect 15106 9560 15162 9616
rect 15106 8880 15162 8936
rect 15106 8200 15162 8256
rect 14462 7520 14518 7576
rect 15106 6840 15162 6896
rect 15198 6196 15200 6216
rect 15200 6196 15252 6216
rect 15252 6196 15254 6216
rect 15198 6160 15254 6196
rect 14462 5480 14518 5536
rect 15106 3476 15108 3496
rect 15108 3476 15160 3496
rect 15160 3476 15162 3496
rect 15106 3440 15162 3476
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 0 15058 800 15088
rect 7373 15058 7439 15061
rect 0 15056 7439 15058
rect 0 15000 7378 15056
rect 7434 15000 7439 15056
rect 0 14998 7439 15000
rect 0 14968 800 14998
rect 7373 14995 7439 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 14825 13018 14891 13021
rect 15806 13018 16606 13048
rect 14825 13016 16606 13018
rect 14825 12960 14830 13016
rect 14886 12960 16606 13016
rect 14825 12958 16606 12960
rect 0 12928 800 12958
rect 14825 12955 14891 12958
rect 15806 12928 16606 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 0 12338 800 12368
rect 15193 12338 15259 12341
rect 15806 12338 16606 12368
rect 0 12248 858 12338
rect 15193 12336 16606 12338
rect 15193 12280 15198 12336
rect 15254 12280 16606 12336
rect 15193 12278 16606 12280
rect 15193 12275 15259 12278
rect 15806 12248 16606 12278
rect 798 12205 858 12248
rect 798 12200 907 12205
rect 798 12144 846 12200
rect 902 12144 907 12200
rect 798 12142 907 12144
rect 841 12139 907 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 841 11794 907 11797
rect 798 11792 907 11794
rect 798 11736 846 11792
rect 902 11736 907 11792
rect 798 11731 907 11736
rect 798 11688 858 11731
rect 0 11598 858 11688
rect 15101 11658 15167 11661
rect 15806 11658 16606 11688
rect 15101 11656 16606 11658
rect 15101 11600 15106 11656
rect 15162 11600 16606 11656
rect 15101 11598 16606 11600
rect 0 11568 800 11598
rect 15101 11595 15167 11598
rect 15806 11568 16606 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 2221 11250 2287 11253
rect 4337 11250 4403 11253
rect 6453 11250 6519 11253
rect 2221 11248 6519 11250
rect 2221 11192 2226 11248
rect 2282 11192 4342 11248
rect 4398 11192 6458 11248
rect 6514 11192 6519 11248
rect 2221 11190 6519 11192
rect 2221 11187 2287 11190
rect 4337 11187 4403 11190
rect 6453 11187 6519 11190
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 15193 10978 15259 10981
rect 15806 10978 16606 11008
rect 15193 10976 16606 10978
rect 15193 10920 15198 10976
rect 15254 10920 16606 10976
rect 15193 10918 16606 10920
rect 15193 10915 15259 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 15806 10888 16606 10918
rect 4870 10847 5186 10848
rect 841 10434 907 10437
rect 798 10432 907 10434
rect 798 10376 846 10432
rect 902 10376 907 10432
rect 798 10371 907 10376
rect 798 10328 858 10371
rect 0 10238 858 10328
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 15101 10298 15167 10301
rect 15806 10298 16606 10328
rect 15101 10296 16606 10298
rect 15101 10240 15106 10296
rect 15162 10240 16606 10296
rect 15101 10238 16606 10240
rect 0 10208 800 10238
rect 15101 10235 15167 10238
rect 15806 10208 16606 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 2221 9618 2287 9621
rect 0 9616 2287 9618
rect 0 9560 2226 9616
rect 2282 9560 2287 9616
rect 0 9558 2287 9560
rect 0 9528 800 9558
rect 2221 9555 2287 9558
rect 15101 9618 15167 9621
rect 15806 9618 16606 9648
rect 15101 9616 16606 9618
rect 15101 9560 15106 9616
rect 15162 9560 16606 9616
rect 15101 9558 16606 9560
rect 15101 9555 15167 9558
rect 15806 9528 16606 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 15101 8938 15167 8941
rect 15806 8938 16606 8968
rect 15101 8936 16606 8938
rect 15101 8880 15106 8936
rect 15162 8880 16606 8936
rect 15101 8878 16606 8880
rect 0 8848 800 8878
rect 15101 8875 15167 8878
rect 15806 8848 16606 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8258 800 8288
rect 1393 8258 1459 8261
rect 0 8256 1459 8258
rect 0 8200 1398 8256
rect 1454 8200 1459 8256
rect 0 8198 1459 8200
rect 0 8168 800 8198
rect 1393 8195 1459 8198
rect 15101 8258 15167 8261
rect 15806 8258 16606 8288
rect 15101 8256 16606 8258
rect 15101 8200 15106 8256
rect 15162 8200 16606 8256
rect 15101 8198 16606 8200
rect 15101 8195 15167 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 15806 8168 16606 8198
rect 4210 8127 4526 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 14457 7578 14523 7581
rect 15806 7578 16606 7608
rect 14457 7576 16606 7578
rect 14457 7520 14462 7576
rect 14518 7520 16606 7576
rect 14457 7518 16606 7520
rect 0 7488 800 7518
rect 14457 7515 14523 7518
rect 15806 7488 16606 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 15101 6898 15167 6901
rect 15806 6898 16606 6928
rect 15101 6896 16606 6898
rect 15101 6840 15106 6896
rect 15162 6840 16606 6896
rect 15101 6838 16606 6840
rect 15101 6835 15167 6838
rect 15806 6808 16606 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 15193 6218 15259 6221
rect 15806 6218 16606 6248
rect 15193 6216 16606 6218
rect 15193 6160 15198 6216
rect 15254 6160 16606 6216
rect 15193 6158 16606 6160
rect 0 6128 800 6158
rect 15193 6155 15259 6158
rect 15806 6128 16606 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 14457 5538 14523 5541
rect 15806 5538 16606 5568
rect 14457 5536 16606 5538
rect 14457 5480 14462 5536
rect 14518 5480 16606 5536
rect 14457 5478 16606 5480
rect 14457 5475 14523 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 15806 5448 16606 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 15101 3498 15167 3501
rect 15806 3498 16606 3528
rect 15101 3496 16606 3498
rect 15101 3440 15106 3496
rect 15162 3440 16606 3496
rect 15101 3438 16606 3440
rect 15101 3435 15167 3438
rect 15806 3408 16606 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 15808 4528 16368
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 16352 5188 16368
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _236_
timestamp 0
transform -1 0 2300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 0
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _238_
timestamp 0
transform -1 0 4416 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _239_
timestamp 0
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _240_
timestamp 0
transform -1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _241_
timestamp 0
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _242_
timestamp 0
transform -1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _243_
timestamp 0
transform -1 0 14996 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _244_
timestamp 0
transform 1 0 9108 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _245_
timestamp 0
transform 1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _246_
timestamp 0
transform 1 0 8188 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _247_
timestamp 0
transform 1 0 8280 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _248_
timestamp 0
transform -1 0 11224 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _249_
timestamp 0
transform -1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _250_
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _251_
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _252_
timestamp 0
transform -1 0 14720 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _253_
timestamp 0
transform -1 0 14996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _254_
timestamp 0
transform 1 0 14720 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _255_
timestamp 0
transform -1 0 14720 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _256_
timestamp 0
transform -1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _257_
timestamp 0
transform 1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _258_
timestamp 0
transform 1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 0
transform -1 0 14996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 0
transform 1 0 14720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 0
transform -1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 0
transform -1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 0
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 0
transform -1 0 5060 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 0
transform 1 0 2576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 0
transform -1 0 14720 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _267_
timestamp 0
transform -1 0 10120 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _268_
timestamp 0
transform -1 0 10580 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _269_
timestamp 0
transform 1 0 8740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _270_
timestamp 0
transform 1 0 8096 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _271_
timestamp 0
transform 1 0 9292 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _272_
timestamp 0
transform -1 0 10120 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _273_
timestamp 0
transform -1 0 9292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _274_
timestamp 0
transform 1 0 9292 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _275_
timestamp 0
transform 1 0 11868 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _276_
timestamp 0
transform -1 0 11868 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _277_
timestamp 0
transform -1 0 13432 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _278_
timestamp 0
transform 1 0 11500 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _279_
timestamp 0
transform 1 0 14168 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _280_
timestamp 0
transform -1 0 14720 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _281_
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _282_
timestamp 0
transform 1 0 13984 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _283_
timestamp 0
transform -1 0 14720 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _284_
timestamp 0
transform 1 0 13432 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _285_
timestamp 0
transform -1 0 14720 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _286_
timestamp 0
transform 1 0 13800 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _287_
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _288_
timestamp 0
transform -1 0 14720 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _289_
timestamp 0
transform 1 0 13432 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _290_
timestamp 0
transform 1 0 14168 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _291_
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _292_
timestamp 0
transform 1 0 12144 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _293_
timestamp 0
transform -1 0 11224 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _294_
timestamp 0
transform 1 0 10488 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _295_
timestamp 0
transform 1 0 8188 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _296_
timestamp 0
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _297_
timestamp 0
transform -1 0 9384 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _298_
timestamp 0
transform 1 0 8004 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _299_
timestamp 0
transform -1 0 10304 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _300_
timestamp 0
transform -1 0 9568 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _301_
timestamp 0
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _302_
timestamp 0
transform 1 0 2576 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _303_
timestamp 0
transform 1 0 4508 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _304_
timestamp 0
transform 1 0 3956 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _305_
timestamp 0
transform -1 0 5060 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _306_
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _307_
timestamp 0
transform 1 0 1748 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _308_
timestamp 0
transform 1 0 1472 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _309_
timestamp 0
transform 1 0 3128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _310_
timestamp 0
transform -1 0 2300 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _311_
timestamp 0
transform 1 0 1472 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _312_
timestamp 0
transform 1 0 2208 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _313_
timestamp 0
transform 1 0 2116 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _314_
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _315_
timestamp 0
transform 1 0 2024 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _316_
timestamp 0
transform 1 0 2668 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _317_
timestamp 0
transform 1 0 3312 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _318_
timestamp 0
transform 1 0 1748 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _319_
timestamp 0
transform 1 0 1472 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _320_
timestamp 0
transform 1 0 3220 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _321_
timestamp 0
transform 1 0 1656 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _322_
timestamp 0
transform 1 0 2024 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _323_
timestamp 0
transform -1 0 3588 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _324_
timestamp 0
transform 1 0 2300 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _325_
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _326_
timestamp 0
transform 1 0 2760 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _327_
timestamp 0
transform -1 0 4324 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _328_
timestamp 0
transform 1 0 3772 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _329_
timestamp 0
transform -1 0 2116 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _330_
timestamp 0
transform 1 0 3864 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _331_
timestamp 0
transform 1 0 3036 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_4  _332_
timestamp 0
transform 1 0 2760 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__or4_4  _333_
timestamp 0
transform 1 0 2852 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _334_
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _335_
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _336_
timestamp 0
transform -1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _337_
timestamp 0
transform -1 0 8096 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _338_
timestamp 0
transform -1 0 3036 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _339_
timestamp 0
transform -1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _340_
timestamp 0
transform -1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _341_
timestamp 0
transform 1 0 3220 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _342_
timestamp 0
transform 1 0 3680 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _343_
timestamp 0
transform 1 0 7728 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _344_
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _345_
timestamp 0
transform -1 0 2576 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _346_
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _347_
timestamp 0
transform 1 0 12420 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _348_
timestamp 0
transform 1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _349_
timestamp 0
transform 1 0 12512 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _350_
timestamp 0
transform 1 0 12144 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _351_
timestamp 0
transform 1 0 12144 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _352_
timestamp 0
transform 1 0 11684 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _353_
timestamp 0
transform 1 0 12696 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _354_
timestamp 0
transform -1 0 13984 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _355_
timestamp 0
transform -1 0 12696 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _356_
timestamp 0
transform 1 0 10856 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _357_
timestamp 0
transform 1 0 10948 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _358_
timestamp 0
transform -1 0 11960 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _359_
timestamp 0
transform -1 0 12144 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _360_
timestamp 0
transform -1 0 12696 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _361_
timestamp 0
transform -1 0 12788 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _362_
timestamp 0
transform 1 0 11592 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _363_
timestamp 0
transform -1 0 11316 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _364_
timestamp 0
transform -1 0 10764 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _365_
timestamp 0
transform -1 0 10212 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _366_
timestamp 0
transform 1 0 11684 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _367_
timestamp 0
transform -1 0 12328 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _368_
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _369_
timestamp 0
transform 1 0 12328 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _370_
timestamp 0
transform 1 0 12788 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _371_
timestamp 0
transform 1 0 12512 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _372_
timestamp 0
transform 1 0 12788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _373_
timestamp 0
transform -1 0 13984 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _374_
timestamp 0
transform 1 0 11592 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _375_
timestamp 0
transform 1 0 12144 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _376_
timestamp 0
transform -1 0 12052 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _377_
timestamp 0
transform -1 0 12512 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _378_
timestamp 0
transform -1 0 10856 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _379_
timestamp 0
transform -1 0 11316 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _380_
timestamp 0
transform -1 0 12144 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _381_
timestamp 0
transform 1 0 9476 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _382_
timestamp 0
transform -1 0 7912 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _383_
timestamp 0
transform -1 0 8096 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _384_
timestamp 0
transform 1 0 7084 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _385_
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _386_
timestamp 0
transform -1 0 8372 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _387_
timestamp 0
transform -1 0 7452 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _388_
timestamp 0
transform -1 0 6808 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _389_
timestamp 0
transform -1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _390_
timestamp 0
transform -1 0 5980 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _391_
timestamp 0
transform -1 0 9016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and4_2  _392_
timestamp 0
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _393_
timestamp 0
transform 1 0 6900 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _394_
timestamp 0
transform 1 0 6808 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _395_
timestamp 0
transform 1 0 9108 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _396_
timestamp 0
transform 1 0 9292 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _397_
timestamp 0
transform 1 0 9568 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _398_
timestamp 0
transform -1 0 9568 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _399_
timestamp 0
transform 1 0 10212 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _400_
timestamp 0
transform 1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _401_
timestamp 0
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _402_
timestamp 0
transform -1 0 8832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _403_
timestamp 0
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _404_
timestamp 0
transform 1 0 8464 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _405_
timestamp 0
transform -1 0 6072 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _406_
timestamp 0
transform 1 0 5520 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _407_
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _408_
timestamp 0
transform -1 0 5520 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _409_
timestamp 0
transform 1 0 5336 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _410_
timestamp 0
transform -1 0 4784 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _411_
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _412_
timestamp 0
transform 1 0 3312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _413_
timestamp 0
transform 1 0 4600 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _414_
timestamp 0
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _415_
timestamp 0
transform -1 0 3220 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _416_
timestamp 0
transform 1 0 5336 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _417_
timestamp 0
transform -1 0 5980 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _418_
timestamp 0
transform 1 0 5060 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _419_
timestamp 0
transform 1 0 5244 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _420_
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _421_
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _422_
timestamp 0
transform 1 0 5336 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _423_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _424_
timestamp 0
transform -1 0 6256 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _425_
timestamp 0
transform -1 0 7360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _426_
timestamp 0
transform -1 0 6992 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _427_
timestamp 0
transform 1 0 4784 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _428_
timestamp 0
transform 1 0 4600 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _429_
timestamp 0
transform -1 0 5244 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _430_
timestamp 0
transform 1 0 4140 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _431_
timestamp 0
transform -1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _432_
timestamp 0
transform -1 0 5060 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _433_
timestamp 0
transform -1 0 4784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _434_
timestamp 0
transform -1 0 4416 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _435_
timestamp 0
transform 1 0 3864 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _436_
timestamp 0
transform -1 0 4232 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _437_
timestamp 0
transform 1 0 4232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _438_
timestamp 0
transform -1 0 4232 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _439_
timestamp 0
transform 1 0 2208 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _440_
timestamp 0
transform 1 0 14904 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _441_
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _442_
timestamp 0
transform -1 0 13800 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _443_
timestamp 0
transform 1 0 10580 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _444_
timestamp 0
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _445_
timestamp 0
transform -1 0 10488 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _446_
timestamp 0
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _447_
timestamp 0
transform -1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 0
transform 1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 0
transform 1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 0
transform -1 0 11592 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 0
transform -1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 0
transform 1 0 7268 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _453_
timestamp 0
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 0
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 0
transform -1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 0
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _457_
timestamp 0
transform -1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _458_
timestamp 0
transform 1 0 7176 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _459_
timestamp 0
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 0
transform -1 0 5888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _461_
timestamp 0
transform -1 0 3680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _462_
timestamp 0
transform 1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _463_
timestamp 0
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _464_
timestamp 0
transform -1 0 7636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _465_
timestamp 0
transform -1 0 9476 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 0
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 0
transform -1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 0
transform -1 0 7452 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 0
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 0
transform -1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _471_
timestamp 0
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _472_
timestamp 0
transform 1 0 12512 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _473_
timestamp 0
transform 1 0 12972 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _474_
timestamp 0
transform 1 0 12144 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _475_
timestamp 0
transform 1 0 11684 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _476_
timestamp 0
transform 1 0 9568 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _477_
timestamp 0
transform 1 0 12144 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _478_
timestamp 0
transform 1 0 9016 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _479_
timestamp 0
transform 1 0 12144 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _480_
timestamp 0
transform 1 0 12144 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _481_
timestamp 0
transform 1 0 12696 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _482_
timestamp 0
transform 1 0 9476 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _483_
timestamp 0
transform 1 0 9476 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _484_
timestamp 0
transform -1 0 9568 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _485_
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _486_
timestamp 0
transform 1 0 5244 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _487_
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _488_
timestamp 0
transform -1 0 11408 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _489_
timestamp 0
transform 1 0 9568 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _490_
timestamp 0
transform 1 0 8464 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _491_
timestamp 0
transform 1 0 6164 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _492_
timestamp 0
transform -1 0 8188 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _493_
timestamp 0
transform 1 0 3772 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _494_
timestamp 0
transform 1 0 1564 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _495_
timestamp 0
transform -1 0 8188 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _496_
timestamp 0
transform -1 0 8188 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _497_
timestamp 0
transform 1 0 6256 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _498_
timestamp 0
transform 1 0 6992 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _499_
timestamp 0
transform 1 0 4232 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _500_
timestamp 0
transform 1 0 5060 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _501_
timestamp 0
transform 1 0 4416 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _502_
timestamp 0
transform 1 0 3496 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _503_
timestamp 0
transform -1 0 3312 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _504_
timestamp 0
transform 1 0 1932 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 7360 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 8648 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform 1 0 10212 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform -1 0 6900 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 9752 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_2  clkload0
timestamp 0
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload1
timestamp 0
transform 1 0 10212 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload2
timestamp 0
transform 1 0 9384 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clone2
timestamp 0
transform -1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout35
timestamp 0
transform -1 0 6072 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout36
timestamp 0
transform 1 0 10672 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout37
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout38
timestamp 0
transform -1 0 10672 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout39
timestamp 0
transform 1 0 14168 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout40
timestamp 0
transform 1 0 13340 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout41
timestamp 0
transform -1 0 13800 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 0
transform -1 0 13800 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16
timestamp 0
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20
timestamp 0
transform 1 0 2944 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 0
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44
timestamp 0
transform 1 0 5152 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76
timestamp 0
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 0
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 0
transform 1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_82
timestamp 0
transform 1 0 8648 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_94
timestamp 0
transform 1 0 9752 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 0
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_121
timestamp 0
transform 1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_148
timestamp 0
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_152
timestamp 0
transform 1 0 15088 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_40
timestamp 0
transform 1 0 4784 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_127
timestamp 0
transform 1 0 12788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 0
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_23
timestamp 0
transform 1 0 3220 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_30
timestamp 0
transform 1 0 3864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 0
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 0
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_48
timestamp 0
transform 1 0 5520 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 0
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_62
timestamp 0
transform 1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_73
timestamp 0
transform 1 0 7820 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_79
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 0
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_75
timestamp 0
transform 1 0 8004 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_88
timestamp 0
transform 1 0 9200 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_99
timestamp 0
transform 1 0 10212 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_111
timestamp 0
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_128
timestamp 0
transform 1 0 12880 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_148
timestamp 0
transform 1 0 14720 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_152
timestamp 0
transform 1 0 15088 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_61
timestamp 0
transform 1 0 6716 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_65
timestamp 0
transform 1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_79
timestamp 0
transform 1 0 8372 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_116
timestamp 0
transform 1 0 11776 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_126
timestamp 0
transform 1 0 12696 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_132
timestamp 0
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_140
timestamp 0
transform 1 0 13984 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_144
timestamp 0
transform 1 0 14352 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_151
timestamp 0
transform 1 0 14996 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_38
timestamp 0
transform 1 0 4600 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_57
timestamp 0
transform 1 0 6348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 0
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 0
transform 1 0 9384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_104
timestamp 0
transform 1 0 10672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_112
timestamp 0
transform 1 0 11408 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 0
transform 1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_6
timestamp 0
transform 1 0 1656 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_22
timestamp 0
transform 1 0 3128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 0
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 0
transform 1 0 8924 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_116
timestamp 0
transform 1 0 11776 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_124
timestamp 0
transform 1 0 12512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_130
timestamp 0
transform 1 0 13064 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_147
timestamp 0
transform 1 0 14628 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 0
transform 1 0 14996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_13
timestamp 0
transform 1 0 2300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 0
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_32
timestamp 0
transform 1 0 4048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_40
timestamp 0
transform 1 0 4784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_61
timestamp 0
transform 1 0 6716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_73
timestamp 0
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 0
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_94
timestamp 0
transform 1 0 9752 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_98
timestamp 0
transform 1 0 10120 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_148
timestamp 0
transform 1 0 14720 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_22
timestamp 0
transform 1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_33
timestamp 0
transform 1 0 4140 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp 0
transform 1 0 5244 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 0
transform 1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_92
timestamp 0
transform 1 0 9568 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_98
timestamp 0
transform 1 0 10120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_138
timestamp 0
transform 1 0 13800 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_144
timestamp 0
transform 1 0 14352 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 0
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_13
timestamp 0
transform 1 0 2300 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_36
timestamp 0
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_40
timestamp 0
transform 1 0 4784 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 0
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_100
timestamp 0
transform 1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_111
timestamp 0
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_123
timestamp 0
transform 1 0 12420 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_135
timestamp 0
transform 1 0 13524 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_148
timestamp 0
transform 1 0 14720 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_6
timestamp 0
transform 1 0 1656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_13
timestamp 0
transform 1 0 2300 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_36
timestamp 0
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 0
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_60
timestamp 0
transform 1 0 6624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_64
timestamp 0
transform 1 0 6992 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_71
timestamp 0
transform 1 0 7636 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 0
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_118
timestamp 0
transform 1 0 11960 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_130
timestamp 0
transform 1 0 13064 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_6
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_37
timestamp 0
transform 1 0 4508 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_45
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_98
timestamp 0
transform 1 0 10120 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_113
timestamp 0
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_148
timestamp 0
transform 1 0 14720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_10
timestamp 0
transform 1 0 2024 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_25
timestamp 0
transform 1 0 3404 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_13_47
timestamp 0
transform 1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 0
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_91
timestamp 0
transform 1 0 9476 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_104
timestamp 0
transform 1 0 10672 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 0
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_126
timestamp 0
transform 1 0 12696 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_130
timestamp 0
transform 1 0 13064 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_134
timestamp 0
transform 1 0 13432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_142
timestamp 0
transform 1 0 14168 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 0
transform 1 0 14996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_13
timestamp 0
transform 1 0 2300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 0
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 0
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_54
timestamp 0
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_111
timestamp 0
transform 1 0 11316 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_127
timestamp 0
transform 1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 0
transform 1 0 14720 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_6
timestamp 0
transform 1 0 1656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_14
timestamp 0
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_35
timestamp 0
transform 1 0 4324 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_43
timestamp 0
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_60
timestamp 0
transform 1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_66
timestamp 0
transform 1 0 7176 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_78
timestamp 0
transform 1 0 8280 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_90
timestamp 0
transform 1 0 9384 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_140
timestamp 0
transform 1 0 13984 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 0
transform 1 0 14996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 0
transform 1 0 1656 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_10
timestamp 0
transform 1 0 2024 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_63
timestamp 0
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_88
timestamp 0
transform 1 0 9200 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_100
timestamp 0
transform 1 0 10304 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_104
timestamp 0
transform 1 0 10672 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_112
timestamp 0
transform 1 0 11408 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_122
timestamp 0
transform 1 0 12328 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_130
timestamp 0
transform 1 0 13064 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 0
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_144
timestamp 0
transform 1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_6
timestamp 0
transform 1 0 1656 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_28
timestamp 0
transform 1 0 3680 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_61
timestamp 0
transform 1 0 6716 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_90
timestamp 0
transform 1 0 9384 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_129
timestamp 0
transform 1 0 12972 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_140
timestamp 0
transform 1 0 13984 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_144
timestamp 0
transform 1 0 14352 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_151
timestamp 0
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_12
timestamp 0
transform 1 0 2208 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_76
timestamp 0
transform 1 0 8096 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 0
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_119
timestamp 0
transform 1 0 12052 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 0
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_26
timestamp 0
transform 1 0 3496 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_38
timestamp 0
transform 1 0 4600 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_50
timestamp 0
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_19_92
timestamp 0
transform 1 0 9568 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_98
timestamp 0
transform 1 0 10120 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 0
transform 1 0 12144 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_130
timestamp 0
transform 1 0 13064 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_136
timestamp 0
transform 1 0 13616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 0
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_152
timestamp 0
transform 1 0 15088 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_6
timestamp 0
transform 1 0 1656 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_21
timestamp 0
transform 1 0 3036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_40
timestamp 0
transform 1 0 4784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_44
timestamp 0
transform 1 0 5152 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_68
timestamp 0
transform 1 0 7360 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 0
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_20_117
timestamp 0
transform 1 0 11868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_130
timestamp 0
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 0
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 0
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp 0
transform 1 0 5336 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp 0
transform 1 0 8372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 0
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_98
timestamp 0
transform 1 0 10120 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 0
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_152
timestamp 0
transform 1 0 15088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_14
timestamp 0
transform 1 0 2392 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_19
timestamp 0
transform 1 0 2852 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_34
timestamp 0
transform 1 0 4232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_46
timestamp 0
transform 1 0 5336 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_58
timestamp 0
transform 1 0 6440 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_66
timestamp 0
transform 1 0 7176 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_70
timestamp 0
transform 1 0 7544 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 0
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_101
timestamp 0
transform 1 0 10396 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_116
timestamp 0
transform 1 0 11776 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_128
timestamp 0
transform 1 0 12880 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_80
timestamp 0
transform 1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_98
timestamp 0
transform 1 0 10120 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 0
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_134
timestamp 0
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_146
timestamp 0
transform 1 0 14536 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_152
timestamp 0
transform 1 0 15088 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_73
timestamp 0
transform 1 0 7820 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_103
timestamp 0
transform 1 0 10580 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_123
timestamp 0
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 0
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_29
timestamp 0
transform 1 0 3772 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_41
timestamp 0
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 0
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_77
timestamp 0
transform 1 0 8188 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_83
timestamp 0
transform 1 0 8740 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_85
timestamp 0
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_90
timestamp 0
transform 1 0 9384 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_104
timestamp 0
transform 1 0 10672 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_118
timestamp 0
transform 1 0 11960 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_130
timestamp 0
transform 1 0 13064 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 0
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_141
timestamp 0
transform 1 0 14076 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 4508 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 14720 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 11316 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform -1 0 11960 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 8740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform 1 0 9108 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform 1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform 1 0 10120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform 1 0 14904 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 0
transform 1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 0
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 0
transform -1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 0
transform 1 0 14904 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 0
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 0
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform 1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 0
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 0
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 0
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 0
transform 1 0 2024 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 0
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 0
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 0
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 0
transform -1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 0
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 0
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 0
transform -1 0 14720 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 0
transform 1 0 14904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 0
transform 1 0 14904 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 0
transform 1 0 14628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 0
transform 1 0 14904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 0
transform -1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 0
transform -1 0 14904 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 0
transform -1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 0
transform 1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_26
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 15456 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_27
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_28
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_29
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_30
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_31
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_32
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 15456 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_33
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_34
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_35
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_36
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_37
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_38
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 15456 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_39
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 15456 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_40
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 15456 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_41
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 15456 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_42
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 15456 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_43
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_44
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_45
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 0
transform -1 0 15456 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_46
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 0
transform -1 0 15456 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_47
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 0
transform -1 0 15456 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_48
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 0
transform -1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_49
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 0
transform -1 0 15456 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_50
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 0
transform -1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_51
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 0
transform -1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1
timestamp 0
transform 1 0 1748 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 0
transform 1 0 2576 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer4
timestamp 0
transform 1 0 3036 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer5
timestamp 0
transform -1 0 2760 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_52
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_53
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_55
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_57
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_58
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_59
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_60
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_61
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_64
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_65
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_67
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_68
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_69
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_70
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_72
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_73
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_74
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_75
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_76
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_77
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_78
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_79
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_80
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_81
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_82
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_83
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_84
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_85
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_86
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_87
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_88
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_89
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_90
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_91
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_92
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_93
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_94
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_95
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_96
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_97
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_98
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_99
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_100
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_101
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_102
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_103
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_104
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_105
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_106
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_107
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_108
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_109
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_110
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_111
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_112
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_113
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_114
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_115
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_116
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_117
timestamp 0
transform 1 0 3680 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_118
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_119
timestamp 0
transform 1 0 8832 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_120
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_121
timestamp 0
transform 1 0 13984 0 -1 16320
box -38 -48 130 592
<< labels >>
rlabel metal1 s 8280 16320 8280 16320 4 VGND
rlabel metal1 s 8280 15776 8280 15776 4 VPWR
rlabel metal2 s 12834 3162 12834 3162 4 _000_
rlabel metal1 s 10028 12614 10028 12614 4 _001_
rlabel metal2 s 9798 13566 9798 13566 4 _002_
rlabel metal1 s 8464 12750 8464 12750 4 _003_
rlabel metal1 s 6762 14042 6762 14042 4 _004_
rlabel metal2 s 5566 13532 5566 13532 4 _005_
rlabel metal2 s 7314 11356 7314 11356 4 _006_
rlabel metal1 s 10626 5882 10626 5882 4 _007_
rlabel metal1 s 10028 4726 10028 4726 4 _008_
rlabel metal2 s 8786 4318 8786 4318 4 _009_
rlabel metal1 s 6486 4488 6486 4488 4 _010_
rlabel metal1 s 13110 4046 13110 4046 4 _011_
rlabel metal2 s 7866 3230 7866 3230 4 _012_
rlabel metal2 s 4094 3230 4094 3230 4 _013_
rlabel metal1 s 1886 4488 1886 4488 4 _014_
rlabel metal1 s 6854 6222 6854 6222 4 _015_
rlabel metal2 s 7866 7582 7866 7582 4 _016_
rlabel metal1 s 6394 8874 6394 8874 4 _017_
rlabel metal1 s 7130 9962 7130 9962 4 _018_
rlabel metal1 s 4692 9690 4692 9690 4 _019_
rlabel metal1 s 5198 11050 5198 11050 4 _020_
rlabel metal1 s 4738 11832 4738 11832 4 _021_
rlabel metal1 s 12466 5576 12466 5576 4 _022_
rlabel metal2 s 3818 14110 3818 14110 4 _023_
rlabel metal2 s 2990 13668 2990 13668 4 _024_
rlabel metal1 s 12052 6970 12052 6970 4 _025_
rlabel metal1 s 10718 8398 10718 8398 4 _026_
rlabel metal2 s 12466 9214 12466 9214 4 _027_
rlabel metal2 s 9338 10268 9338 10268 4 _028_
rlabel metal1 s 12098 10540 12098 10540 4 _029_
rlabel metal1 s 12696 11594 12696 11594 4 _030_
rlabel metal2 s 12742 13566 12742 13566 4 _031_
rlabel metal1 s 14313 3094 14313 3094 4 _032_
rlabel metal1 s 15042 4148 15042 4148 4 _033_
rlabel metal2 s 13846 5474 13846 5474 4 _034_
rlabel metal1 s 13439 7446 13439 7446 4 _035_
rlabel metal1 s 10672 8058 10672 8058 4 _036_
rlabel metal1 s 13248 9350 13248 9350 4 _037_
rlabel metal2 s 10350 10200 10350 10200 4 _038_
rlabel metal2 s 14214 10880 14214 10880 4 _039_
rlabel metal2 s 13846 12002 13846 12002 4 _040_
rlabel metal1 s 14451 13974 14451 13974 4 _041_
rlabel metal2 s 10534 11560 10534 11560 4 _042_
rlabel metal1 s 11231 13226 11231 13226 4 _043_
rlabel metal1 s 8648 12410 8648 12410 4 _044_
rlabel metal1 s 7360 14586 7360 14586 4 _045_
rlabel metal2 s 6118 13532 6118 13532 4 _046_
rlabel metal1 s 8793 11050 8793 11050 4 _047_
rlabel metal1 s 11638 6392 11638 6392 4 _048_
rlabel metal1 s 11369 5270 11369 5270 4 _049_
rlabel metal1 s 10173 4114 10173 4114 4 _050_
rlabel metal1 s 7406 4114 7406 4114 4 _051_
rlabel metal2 s 6762 2822 6762 2822 4 _052_
rlabel metal1 s 5527 3094 5527 3094 4 _053_
rlabel metal1 s 3319 4522 3319 4522 4 _054_
rlabel metal1 s 6854 5338 6854 5338 4 _055_
rlabel metal1 s 6854 6834 6854 6834 4 _056_
rlabel metal1 s 7544 8602 7544 8602 4 _057_
rlabel metal2 s 9338 9792 9338 9792 4 _058_
rlabel metal1 s 5336 10438 5336 10438 4 _059_
rlabel metal2 s 6486 10948 6486 10948 4 _060_
rlabel metal2 s 7314 11934 7314 11934 4 _061_
rlabel metal1 s 4738 13498 4738 13498 4 _062_
rlabel metal2 s 2898 13702 2898 13702 4 _063_
rlabel metal1 s 3220 2618 3220 2618 4 _064_
rlabel metal1 s 2162 2618 2162 2618 4 _065_
rlabel metal1 s 1518 7412 1518 7412 4 _066_
rlabel metal1 s 4876 2618 4876 2618 4 _067_
rlabel metal2 s 4278 4318 4278 4318 4 _068_
rlabel metal1 s 3956 6970 3956 6970 4 _069_
rlabel metal2 s 8234 5746 8234 5746 4 _070_
rlabel metal1 s 8832 5610 8832 5610 4 _071_
rlabel metal2 s 9982 7956 9982 7956 4 _072_
rlabel metal1 s 10386 7854 10386 7854 4 _073_
rlabel metal1 s 9936 15538 9936 15538 4 _074_
rlabel metal1 s 9064 14994 9064 14994 4 _075_
rlabel metal1 s 8694 15062 8694 15062 4 _076_
rlabel metal2 s 8326 15028 8326 15028 4 _077_
rlabel metal1 s 11224 15538 11224 15538 4 _078_
rlabel metal1 s 12926 14892 12926 14892 4 _079_
rlabel metal1 s 13156 13294 13156 13294 4 _080_
rlabel metal1 s 14398 12784 14398 12784 4 _081_
rlabel metal2 s 14582 12036 14582 12036 4 _082_
rlabel metal1 s 14628 11526 14628 11526 4 _083_
rlabel metal1 s 14674 10710 14674 10710 4 _084_
rlabel metal1 s 14444 9690 14444 9690 4 _085_
rlabel metal1 s 14582 8602 14582 8602 4 _086_
rlabel metal1 s 14628 7174 14628 7174 4 _087_
rlabel metal2 s 14582 6086 14582 6086 4 _088_
rlabel metal1 s 14214 6324 14214 6324 4 _089_
rlabel metal1 s 14720 5338 14720 5338 4 _090_
rlabel metal2 s 1886 7548 1886 7548 4 _091_
rlabel metal1 s 6762 10030 6762 10030 4 _092_
rlabel metal1 s 3082 11084 3082 11084 4 _093_
rlabel metal2 s 3450 11662 3450 11662 4 _094_
rlabel metal2 s 2622 13770 2622 13770 4 _095_
rlabel metal1 s 9890 15878 9890 15878 4 _096_
rlabel metal1 s 10212 15130 10212 15130 4 _097_
rlabel metal1 s 9430 14994 9430 14994 4 _098_
rlabel metal1 s 9338 15470 9338 15470 4 _099_
rlabel metal1 s 9752 14994 9752 14994 4 _100_
rlabel metal1 s 11086 14416 11086 14416 4 _101_
rlabel metal1 s 9706 15538 9706 15538 4 _102_
rlabel metal1 s 10350 14858 10350 14858 4 _103_
rlabel metal2 s 12742 15164 12742 15164 4 _104_
rlabel metal1 s 11776 15130 11776 15130 4 _105_
rlabel metal2 s 11822 14722 11822 14722 4 _106_
rlabel metal1 s 11822 14586 11822 14586 4 _107_
rlabel metal2 s 14214 14008 14214 14008 4 _108_
rlabel metal2 s 14030 8636 14030 8636 4 _109_
rlabel metal1 s 13984 5882 13984 5882 4 _110_
rlabel metal1 s 13984 6290 13984 6290 4 _111_
rlabel metal1 s 13662 6324 13662 6324 4 _112_
rlabel metal1 s 13846 6426 13846 6426 4 _113_
rlabel metal1 s 14490 8058 14490 8058 4 _114_
rlabel metal2 s 13846 9248 13846 9248 4 _115_
rlabel metal1 s 14030 10030 14030 10030 4 _116_
rlabel metal1 s 13662 10064 13662 10064 4 _117_
rlabel metal2 s 13478 12240 13478 12240 4 _118_
rlabel metal1 s 14766 12410 14766 12410 4 _119_
rlabel metal2 s 10718 14722 10718 14722 4 _120_
rlabel metal1 s 11638 14926 11638 14926 4 _121_
rlabel metal2 s 10994 14586 10994 14586 4 _122_
rlabel metal1 s 10120 14246 10120 14246 4 _123_
rlabel metal1 s 8142 6902 8142 6902 4 _124_
rlabel metal1 s 8372 6970 8372 6970 4 _125_
rlabel metal1 s 8694 5882 8694 5882 4 _126_
rlabel metal2 s 8510 7174 8510 7174 4 _127_
rlabel metal1 s 9338 7854 9338 7854 4 _128_
rlabel metal2 s 9154 7616 9154 7616 4 _129_
rlabel metal1 s 8832 7786 8832 7786 4 _130_
rlabel metal1 s 3680 5814 3680 5814 4 _131_
rlabel metal1 s 4232 6290 4232 6290 4 _132_
rlabel metal1 s 4416 5882 4416 5882 4 _133_
rlabel metal1 s 4646 4794 4646 4794 4 _134_
rlabel metal1 s 3726 7378 3726 7378 4 _135_
rlabel metal2 s 2530 9350 2530 9350 4 _136_
rlabel metal1 s 2116 9350 2116 9350 4 _137_
rlabel metal2 s 3174 9180 3174 9180 4 _138_
rlabel metal2 s 2346 8772 2346 8772 4 _139_
rlabel metal1 s 2254 9520 2254 9520 4 _140_
rlabel metal1 s 3312 8398 3312 8398 4 _141_
rlabel metal2 s 2898 7854 2898 7854 4 _142_
rlabel metal1 s 2925 8398 2925 8398 4 _143_
rlabel metal1 s 2622 6426 2622 6426 4 _144_
rlabel metal1 s 3220 7378 3220 7378 4 _145_
rlabel metal2 s 3726 7684 3726 7684 4 _146_
rlabel metal1 s 3174 12750 3174 12750 4 _147_
rlabel metal1 s 2530 12750 2530 12750 4 _148_
rlabel metal1 s 2530 11764 2530 11764 4 _149_
rlabel metal2 s 2323 12342 2323 12342 4 _150_
rlabel metal1 s 2622 12614 2622 12614 4 _151_
rlabel metal2 s 2806 11900 2806 11900 4 _152_
rlabel metal1 s 2714 11220 2714 11220 4 _153_
rlabel metal2 s 4738 9418 4738 9418 4 _154_
rlabel metal1 s 3036 10574 3036 10574 4 _155_
rlabel metal2 s 3818 8942 3818 8942 4 _156_
rlabel metal1 s 3542 7242 3542 7242 4 _157_
rlabel metal2 s 2070 7650 2070 7650 4 _158_
rlabel metal1 s 3634 6290 3634 6290 4 _159_
rlabel metal1 s 3910 7718 3910 7718 4 _160_
rlabel metal2 s 3082 10030 3082 10030 4 _161_
rlabel metal1 s 3680 8398 3680 8398 4 _162_
rlabel metal1 s 8050 7956 8050 7956 4 _163_
rlabel metal1 s 9706 8058 9706 8058 4 _164_
rlabel metal1 s 8418 7514 8418 7514 4 _165_
rlabel metal1 s 7728 8058 7728 8058 4 _166_
rlabel metal2 s 2990 9248 2990 9248 4 _167_
rlabel metal2 s 2806 10506 2806 10506 4 _168_
rlabel metal1 s 3128 9690 3128 9690 4 _169_
rlabel metal1 s 3956 6426 3956 6426 4 _170_
rlabel metal1 s 8050 8432 8050 8432 4 _171_
rlabel metal2 s 8510 8738 8510 8738 4 _172_
rlabel metal2 s 6486 9843 6486 9843 4 _173_
rlabel metal2 s 12742 4182 12742 4182 4 _174_
rlabel metal1 s 12612 4250 12612 4250 4 _175_
rlabel metal1 s 12052 5338 12052 5338 4 _176_
rlabel metal1 s 11976 5610 11976 5610 4 _177_
rlabel metal1 s 12512 6630 12512 6630 4 _178_
rlabel metal1 s 13018 6834 13018 6834 4 _179_
rlabel metal1 s 11362 8058 11362 8058 4 _180_
rlabel metal1 s 11625 8602 11625 8602 4 _181_
rlabel metal2 s 12098 9248 12098 9248 4 _182_
rlabel metal1 s 12558 9962 12558 9962 4 _183_
rlabel metal2 s 11270 10336 11270 10336 4 _184_
rlabel metal1 s 10442 10234 10442 10234 4 _185_
rlabel metal1 s 10250 10778 10250 10778 4 _186_
rlabel metal2 s 11914 10710 11914 10710 4 _187_
rlabel metal1 s 11776 12954 11776 12954 4 _188_
rlabel metal2 s 12742 12070 12742 12070 4 _189_
rlabel metal1 s 12880 13294 12880 13294 4 _190_
rlabel metal1 s 12742 13498 12742 13498 4 _191_
rlabel metal1 s 11730 12784 11730 12784 4 _192_
rlabel metal1 s 12098 13294 12098 13294 4 _193_
rlabel metal1 s 11040 12750 11040 12750 4 _194_
rlabel metal1 s 11684 12886 11684 12886 4 _195_
rlabel metal1 s 10396 12954 10396 12954 4 _196_
rlabel metal1 s 9844 13838 9844 13838 4 _197_
rlabel metal2 s 7498 13702 7498 13702 4 _198_
rlabel metal1 s 7590 12410 7590 12410 4 _199_
rlabel metal1 s 7452 13974 7452 13974 4 _200_
rlabel metal1 s 7682 13770 7682 13770 4 _201_
rlabel metal1 s 6072 13702 6072 13702 4 _202_
rlabel metal1 s 7084 13498 7084 13498 4 _203_
rlabel metal1 s 8740 13294 8740 13294 4 _204_
rlabel metal1 s 7774 11730 7774 11730 4 _205_
rlabel metal2 s 7222 11968 7222 11968 4 _206_
rlabel metal1 s 9752 5610 9752 5610 4 _207_
rlabel metal1 s 9660 5814 9660 5814 4 _208_
rlabel metal1 s 9104 4590 9104 4590 4 _209_
rlabel metal1 s 10304 4794 10304 4794 4 _210_
rlabel metal1 s 8280 4590 8280 4590 4 _211_
rlabel metal1 s 6762 4250 6762 4250 4 _212_
rlabel metal1 s 5842 4080 5842 4080 4 _213_
rlabel metal1 s 5612 4250 5612 4250 4 _214_
rlabel metal2 s 5750 3672 5750 3672 4 _215_
rlabel metal2 s 5382 4182 5382 4182 4 _216_
rlabel metal1 s 4278 3536 4278 3536 4 _217_
rlabel metal1 s 3174 3910 3174 3910 4 _218_
rlabel metal1 s 5566 5780 5566 5780 4 _219_
rlabel metal1 s 4178 4250 4178 4250 4 _220_
rlabel metal1 s 5520 5882 5520 5882 4 _221_
rlabel metal1 s 5068 7786 5068 7786 4 _222_
rlabel metal1 s 5428 6970 5428 6970 4 _223_
rlabel metal2 s 5750 7616 5750 7616 4 _224_
rlabel metal1 s 5842 8976 5842 8976 4 _225_
rlabel metal1 s 6900 8534 6900 8534 4 _226_
rlabel metal2 s 7130 9248 7130 9248 4 _227_
rlabel metal1 s 4830 9656 4830 9656 4 _228_
rlabel metal1 s 5144 8602 5144 8602 4 _229_
rlabel metal1 s 4416 9418 4416 9418 4 _230_
rlabel metal1 s 4554 11152 4554 11152 4 _231_
rlabel metal1 s 4416 12138 4416 12138 4 _232_
rlabel metal2 s 3910 12070 3910 12070 4 _233_
rlabel metal1 s 3910 13498 3910 13498 4 _234_
rlabel metal1 s 3542 13158 3542 13158 4 _235_
rlabel metal3 s 4040 15028 4040 15028 4 clk
rlabel metal1 s 9338 12138 9338 12138 4 clknet_0_clk
rlabel metal1 s 1794 3026 1794 3026 4 clknet_2_0__leaf_clk
rlabel metal2 s 13018 4930 13018 4930 4 clknet_2_1__leaf_clk
rlabel metal2 s 5290 14144 5290 14144 4 clknet_2_2__leaf_clk
rlabel metal2 s 9522 13022 9522 13022 4 clknet_2_3__leaf_clk
rlabel metal1 s 14720 5202 14720 5202 4 net1
rlabel metal1 s 8464 2618 8464 2618 4 net10
rlabel metal1 s 8096 2618 8096 2618 4 net11
rlabel metal2 s 14950 6460 14950 6460 4 net12
rlabel metal1 s 1610 10744 1610 10744 4 net13
rlabel metal1 s 5244 4658 5244 4658 4 net14
rlabel metal1 s 5106 2448 5106 2448 4 net15
rlabel metal1 s 1978 6154 1978 6154 4 net16
rlabel metal1 s 1656 7242 1656 7242 4 net17
rlabel metal1 s 1702 7378 1702 7378 4 net18
rlabel metal2 s 1794 9962 1794 9962 4 net19
rlabel metal2 s 13018 15232 13018 15232 4 net2
rlabel metal1 s 1794 8840 1794 8840 4 net20
rlabel metal1 s 1610 11186 1610 11186 4 net21
rlabel metal2 s 2346 11424 2346 11424 4 net22
rlabel metal2 s 14766 5916 14766 5916 4 net23
rlabel metal2 s 1518 13022 1518 13022 4 net24
rlabel metal2 s 1794 12342 1794 12342 4 net25
rlabel metal1 s 14720 7378 14720 7378 4 net26
rlabel metal1 s 14858 8058 14858 8058 4 net27
rlabel metal1 s 14812 9146 14812 9146 4 net28
rlabel metal2 s 14766 10812 14766 10812 4 net29
rlabel metal1 s 12190 15572 12190 15572 4 net3
rlabel metal2 s 14950 11526 14950 11526 4 net30
rlabel metal1 s 14490 12852 14490 12852 4 net31
rlabel metal2 s 14674 14212 14674 14212 4 net32
rlabel metal1 s 13708 8466 13708 8466 4 net33
rlabel metal1 s 4554 2482 4554 2482 4 net34
rlabel metal1 s 2668 2550 2668 2550 4 net35
rlabel metal1 s 9890 4522 9890 4522 4 net36
rlabel metal1 s 4462 14314 4462 14314 4 net37
rlabel metal2 s 12558 11288 12558 11288 4 net38
rlabel metal1 s 3450 2414 3450 2414 4 net39
rlabel metal2 s 8418 15674 8418 15674 4 net4
rlabel metal1 s 13662 5202 13662 5202 4 net40
rlabel metal1 s 13340 9554 13340 9554 4 net41
rlabel metal1 s 14122 13838 14122 13838 4 net42
rlabel metal1 s 2438 14382 2438 14382 4 net43
rlabel metal2 s 4370 11169 4370 11169 4 net44
rlabel metal1 s 3174 12818 3174 12818 4 net45
rlabel metal1 s 3128 11594 3128 11594 4 net46
rlabel metal2 s 2530 10812 2530 10812 4 net47
rlabel metal1 s 8740 15470 8740 15470 4 net5
rlabel metal1 s 2346 2448 2346 2448 4 net59
rlabel metal2 s 10350 15232 10350 15232 4 net6
rlabel metal1 s 10074 15980 10074 15980 4 net7
rlabel metal2 s 14950 9724 14950 9724 4 net8
rlabel metal1 s 14904 8466 14904 8466 4 net9
rlabel metal2 s 3910 1520 3910 1520 4 out
rlabel metal2 s 14490 5355 14490 5355 4 psc[0]
rlabel metal1 s 11040 16082 11040 16082 4 psc[10]
rlabel metal1 s 11684 16082 11684 16082 4 psc[11]
rlabel metal1 s 8464 16082 8464 16082 4 psc[12]
rlabel metal1 s 9200 16082 9200 16082 4 psc[13]
rlabel metal1 s 10534 16082 10534 16082 4 psc[14]
rlabel metal1 s 10350 16116 10350 16116 4 psc[15]
rlabel metal2 s 15134 10149 15134 10149 4 psc[16]
rlabel metal2 s 15134 8687 15134 8687 4 psc[17]
rlabel metal2 s 8418 1588 8418 1588 4 psc[18]
rlabel metal2 s 7774 1588 7774 1588 4 psc[19]
rlabel metal2 s 15134 6817 15134 6817 4 psc[1]
rlabel metal3 s 0 10208 800 10328 4 psc[20]
port 17 nsew
rlabel metal2 s 6486 1554 6486 1554 4 psc[21]
rlabel metal2 s 7130 1027 7130 1027 4 psc[22]
rlabel metal3 s 0 6128 800 6248 4 psc[23]
port 20 nsew
rlabel metal3 s 1050 8228 1050 8228 4 psc[24]
rlabel metal3 s 0 7488 800 7608 4 psc[25]
port 22 nsew
rlabel metal3 s 1464 9588 1464 9588 4 psc[26]
rlabel metal3 s 0 8848 800 8968 4 psc[27]
port 24 nsew
rlabel metal3 s 1050 10948 1050 10948 4 psc[28]
rlabel metal3 s 0 11568 800 11688 4 psc[29]
port 26 nsew
rlabel metal1 s 13202 6256 13202 6256 4 psc[2]
rlabel metal3 s 0 12928 800 13048 4 psc[30]
port 28 nsew
rlabel metal3 s 0 12248 800 12368 4 psc[31]
port 29 nsew
rlabel metal2 s 14490 7463 14490 7463 4 psc[3]
rlabel metal2 s 15134 8041 15134 8041 4 psc[4]
rlabel metal1 s 15134 8964 15134 8964 4 psc[5]
rlabel metal1 s 14858 11084 14858 11084 4 psc[6]
rlabel metal2 s 15134 11373 15134 11373 4 psc[7]
rlabel metal1 s 15180 13294 15180 13294 4 psc[8]
rlabel metal2 s 14858 13141 14858 13141 4 psc[9]
rlabel metal2 s 13110 3298 13110 3298 4 psc_cnt\[0\]
rlabel metal1 s 11546 12138 11546 12138 4 psc_cnt\[10\]
rlabel metal1 s 11178 15436 11178 15436 4 psc_cnt\[11\]
rlabel metal2 s 7774 12954 7774 12954 4 psc_cnt\[12\]
rlabel metal1 s 8188 14994 8188 14994 4 psc_cnt\[13\]
rlabel metal1 s 7314 13430 7314 13430 4 psc_cnt\[14\]
rlabel metal2 s 8786 11526 8786 11526 4 psc_cnt\[15\]
rlabel metal2 s 8786 7956 8786 7956 4 psc_cnt\[16\]
rlabel metal1 s 10488 5610 10488 5610 4 psc_cnt\[17\]
rlabel metal2 s 8970 4250 8970 4250 4 psc_cnt\[18\]
rlabel metal2 s 8326 4998 8326 4998 4 psc_cnt\[19\]
rlabel metal1 s 14030 5678 14030 5678 4 psc_cnt\[1\]
rlabel metal2 s 4278 6460 4278 6460 4 psc_cnt\[20\]
rlabel metal2 s 4554 3230 4554 3230 4 psc_cnt\[21\]
rlabel metal1 s 4784 5678 4784 5678 4 psc_cnt\[22\]
rlabel metal1 s 2530 6188 2530 6188 4 psc_cnt\[23\]
rlabel metal1 s 2208 7310 2208 7310 4 psc_cnt\[24\]
rlabel metal2 s 1978 7344 1978 7344 4 psc_cnt\[25\]
rlabel metal1 s 1794 9554 1794 9554 4 psc_cnt\[26\]
rlabel metal1 s 5842 10166 5842 10166 4 psc_cnt\[27\]
rlabel metal1 s 4830 11118 4830 11118 4 psc_cnt\[28\]
rlabel metal1 s 5612 12206 5612 12206 4 psc_cnt\[29\]
rlabel metal2 s 12466 5746 12466 5746 4 psc_cnt\[2\]
rlabel metal1 s 4462 13328 4462 13328 4 psc_cnt\[30\]
rlabel metal1 s 1610 13838 1610 13838 4 psc_cnt\[31\]
rlabel metal1 s 13846 6766 13846 6766 4 psc_cnt\[3\]
rlabel metal2 s 14490 8432 14490 8432 4 psc_cnt\[4\]
rlabel metal1 s 14260 8942 14260 8942 4 psc_cnt\[5\]
rlabel metal1 s 14628 10234 14628 10234 4 psc_cnt\[6\]
rlabel metal2 s 14306 11390 14306 11390 4 psc_cnt\[7\]
rlabel metal1 s 13018 12852 13018 12852 4 psc_cnt\[8\]
rlabel metal1 s 14858 13872 14858 13872 4 psc_cnt\[9\]
rlabel metal3 s 15134 3485 15134 3485 4 rst
flabel metal4 s 4868 2128 5188 16368 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4208 2128 4528 16368 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 14968 800 15088 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 out
port 4 nsew
flabel metal3 s 15806 5448 16606 5568 0 FreeSans 600 0 0 0 psc[0]
port 5 nsew
flabel metal2 s 10966 17950 11022 18750 0 FreeSans 280 90 0 0 psc[10]
port 6 nsew
flabel metal2 s 11610 17950 11666 18750 0 FreeSans 280 90 0 0 psc[11]
port 7 nsew
flabel metal2 s 8390 17950 8446 18750 0 FreeSans 280 90 0 0 psc[12]
port 8 nsew
flabel metal2 s 9034 17950 9090 18750 0 FreeSans 280 90 0 0 psc[13]
port 9 nsew
flabel metal2 s 10322 17950 10378 18750 0 FreeSans 280 90 0 0 psc[14]
port 10 nsew
flabel metal2 s 9678 17950 9734 18750 0 FreeSans 280 90 0 0 psc[15]
port 11 nsew
flabel metal3 s 15806 10208 16606 10328 0 FreeSans 600 0 0 0 psc[16]
port 12 nsew
flabel metal3 s 15806 8848 16606 8968 0 FreeSans 600 0 0 0 psc[17]
port 13 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 psc[18]
port 14 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 psc[19]
port 15 nsew
flabel metal3 s 15806 6808 16606 6928 0 FreeSans 600 0 0 0 psc[1]
port 16 nsew
flabel metal3 s 400 10268 400 10268 0 FreeSans 600 0 0 0 psc[20]
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 psc[21]
port 18 nsew
flabel metal2 s 7102 0 7158 800 0 FreeSans 280 90 0 0 psc[22]
port 19 nsew
flabel metal3 s 400 6188 400 6188 0 FreeSans 600 0 0 0 psc[23]
flabel metal3 s 0 8168 800 8288 0 FreeSans 600 0 0 0 psc[24]
port 21 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 psc[25]
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 psc[26]
port 23 nsew
flabel metal3 s 400 8908 400 8908 0 FreeSans 600 0 0 0 psc[27]
flabel metal3 s 0 10888 800 11008 0 FreeSans 600 0 0 0 psc[28]
port 25 nsew
flabel metal3 s 400 11628 400 11628 0 FreeSans 600 0 0 0 psc[29]
flabel metal3 s 15806 6128 16606 6248 0 FreeSans 600 0 0 0 psc[2]
port 27 nsew
flabel metal3 s 400 12988 400 12988 0 FreeSans 600 0 0 0 psc[30]
flabel metal3 s 400 12308 400 12308 0 FreeSans 600 0 0 0 psc[31]
flabel metal3 s 15806 7488 16606 7608 0 FreeSans 600 0 0 0 psc[3]
port 30 nsew
flabel metal3 s 15806 8168 16606 8288 0 FreeSans 600 0 0 0 psc[4]
port 31 nsew
flabel metal3 s 15806 9528 16606 9648 0 FreeSans 600 0 0 0 psc[5]
port 32 nsew
flabel metal3 s 15806 10888 16606 11008 0 FreeSans 600 0 0 0 psc[6]
port 33 nsew
flabel metal3 s 15806 11568 16606 11688 0 FreeSans 600 0 0 0 psc[7]
port 34 nsew
flabel metal3 s 15806 12248 16606 12368 0 FreeSans 600 0 0 0 psc[8]
port 35 nsew
flabel metal3 s 15806 12928 16606 13048 0 FreeSans 600 0 0 0 psc[9]
port 36 nsew
flabel metal3 s 15806 3408 16606 3528 0 FreeSans 600 0 0 0 rst
port 37 nsew
<< properties >>
string FIXED_BBOX 0 0 16606 18750
<< end >>
