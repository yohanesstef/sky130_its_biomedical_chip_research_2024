magic
tech sky130A
magscale 1 2
timestamp 1729851530
<< error_p >>
rect -32 525 32 531
rect -32 491 -20 525
rect -32 485 32 491
<< nwell >>
rect -130 -578 130 544
<< pmos >>
rect -36 -516 36 444
<< pdiff >>
rect -94 432 -36 444
rect -94 -504 -82 432
rect -48 -504 -36 432
rect -94 -516 -36 -504
rect 36 432 94 444
rect 36 -504 48 432
rect 82 -504 94 432
rect 36 -516 94 -504
<< pdiffc >>
rect -82 -504 -48 432
rect 48 -504 82 432
<< poly >>
rect -36 525 36 541
rect -36 491 -20 525
rect 20 491 36 525
rect -36 444 36 491
rect -36 -542 36 -516
<< polycont >>
rect -20 491 20 525
<< locali >>
rect -36 491 -20 525
rect 20 491 36 525
rect -82 432 -48 448
rect -82 -520 -48 -504
rect 48 432 82 448
rect 48 -520 82 -504
<< viali >>
rect -20 491 20 525
rect -82 -504 -48 432
rect 48 -504 82 432
<< metal1 >>
rect -32 525 32 531
rect -32 491 -20 525
rect 20 491 32 525
rect -32 485 32 491
rect -88 432 -42 444
rect -88 -504 -82 432
rect -48 -504 -42 432
rect -88 -516 -42 -504
rect 42 432 88 444
rect 42 -504 48 432
rect 82 -504 88 432
rect 42 -516 88 -504
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4.8 l 0.36 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
