VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO freq_psc
  CLASS BLOCK ;
  FOREIGN freq_psc ;
  ORIGIN 0.000 0.000 ;
  SIZE 47.425 BY 58.145 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 46.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 46.480 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END clk
  PIN out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END out
  PIN psc[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 54.145 22.910 58.145 ;
    END
  END psc[0]
  PIN psc[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 54.145 19.690 58.145 ;
    END
  END psc[1]
  PIN psc[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 54.145 32.570 58.145 ;
    END
  END psc[2]
  PIN psc[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.425 34.040 47.425 34.640 ;
    END
  END psc[3]
  PIN psc[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.425 30.640 47.425 31.240 ;
    END
  END psc[4]
  PIN psc[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.425 27.240 47.425 27.840 ;
    END
  END psc[5]
  PIN psc[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.425 13.640 47.425 14.240 ;
    END
  END psc[6]
  PIN psc[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.425 17.040 47.425 17.640 ;
    END
  END psc[7]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END rst
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 42.050 46.430 ;
      LAYER li1 ;
        RECT 5.520 10.795 41.860 46.325 ;
      LAYER met1 ;
        RECT 4.210 10.640 41.860 46.480 ;
      LAYER met2 ;
        RECT 4.230 53.865 19.130 54.810 ;
        RECT 19.970 53.865 22.350 54.810 ;
        RECT 23.190 53.865 32.010 54.810 ;
        RECT 32.850 53.865 40.390 54.810 ;
        RECT 4.230 10.695 40.390 53.865 ;
      LAYER met3 ;
        RECT 3.990 35.040 43.425 46.405 ;
        RECT 4.400 33.640 43.025 35.040 ;
        RECT 3.990 31.640 43.425 33.640 ;
        RECT 4.400 30.240 43.025 31.640 ;
        RECT 3.990 28.240 43.425 30.240 ;
        RECT 3.990 26.840 43.025 28.240 ;
        RECT 3.990 18.040 43.425 26.840 ;
        RECT 4.400 16.640 43.025 18.040 ;
        RECT 3.990 14.640 43.425 16.640 ;
        RECT 3.990 13.240 43.025 14.640 ;
        RECT 3.990 10.715 43.425 13.240 ;
  END
END freq_psc
END LIBRARY

