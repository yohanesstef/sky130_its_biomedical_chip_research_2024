magic
tech sky130A
magscale 1 2
timestamp 1729899137
<< viali >>
rect 3893 9061 3927 9095
rect 4628 8925 4662 8959
rect 4721 8925 4755 8959
rect 4997 8925 5031 8959
rect 5273 8925 5307 8959
rect 6561 8925 6595 8959
rect 3341 8857 3375 8891
rect 4261 8857 4295 8891
rect 3801 8789 3835 8823
rect 4353 8789 4387 8823
rect 4813 8789 4847 8823
rect 5089 8789 5123 8823
rect 6745 8789 6779 8823
rect 4353 8517 4387 8551
rect 7205 8517 7239 8551
rect 6653 8449 6687 8483
rect 6746 8449 6780 8483
rect 7113 8449 7147 8483
rect 7389 8449 7423 8483
rect 4445 8381 4479 8415
rect 4721 8381 4755 8415
rect 7021 8313 7055 8347
rect 3065 8245 3099 8279
rect 6193 8245 6227 8279
rect 7389 8245 7423 8279
rect 3433 8041 3467 8075
rect 4721 8041 4755 8075
rect 5733 8041 5767 8075
rect 6009 8041 6043 8075
rect 3893 7973 3927 8007
rect 7481 7973 7515 8007
rect 6653 7905 6687 7939
rect 7113 7905 7147 7939
rect 3157 7837 3191 7871
rect 4077 7837 4111 7871
rect 4353 7815 4387 7849
rect 4997 7837 5031 7871
rect 5181 7837 5215 7871
rect 5825 7837 5859 7871
rect 5917 7837 5951 7871
rect 6745 7837 6779 7871
rect 7205 7837 7239 7871
rect 7481 7837 7515 7871
rect 2881 7769 2915 7803
rect 3617 7769 3651 7803
rect 4261 7769 4295 7803
rect 4689 7769 4723 7803
rect 4905 7769 4939 7803
rect 7297 7769 7331 7803
rect 1409 7701 1443 7735
rect 3249 7701 3283 7735
rect 3417 7701 3451 7735
rect 4537 7701 4571 7735
rect 5089 7701 5123 7735
rect 6469 7701 6503 7735
rect 6929 7701 6963 7735
rect 7021 7701 7055 7735
rect 2237 7497 2271 7531
rect 3065 7497 3099 7531
rect 4445 7497 4479 7531
rect 6837 7497 6871 7531
rect 7297 7497 7331 7531
rect 2881 7429 2915 7463
rect 3893 7429 3927 7463
rect 4721 7429 4755 7463
rect 2329 7361 2363 7395
rect 2697 7361 2731 7395
rect 3801 7361 3835 7395
rect 3985 7361 4019 7395
rect 4077 7361 4111 7395
rect 4231 7361 4265 7395
rect 5089 7361 5123 7395
rect 7051 7361 7085 7395
rect 7205 7361 7239 7395
rect 8033 7361 8067 7395
rect 7757 7293 7791 7327
rect 4537 7225 4571 7259
rect 7481 7225 7515 7259
rect 7849 7225 7883 7259
rect 4721 7157 4755 7191
rect 4261 6953 4295 6987
rect 4445 6885 4479 6919
rect 3157 6817 3191 6851
rect 4537 6817 4571 6851
rect 4813 6817 4847 6851
rect 3341 6749 3375 6783
rect 3433 6749 3467 6783
rect 3893 6749 3927 6783
rect 6653 6749 6687 6783
rect 6745 6749 6779 6783
rect 7481 6749 7515 6783
rect 2881 6681 2915 6715
rect 3617 6681 3651 6715
rect 1409 6613 1443 6647
rect 4261 6613 4295 6647
rect 6285 6613 6319 6647
rect 7389 6613 7423 6647
rect 2789 6409 2823 6443
rect 5641 6409 5675 6443
rect 2329 6341 2363 6375
rect 3065 6341 3099 6375
rect 5073 6341 5107 6375
rect 5273 6341 5307 6375
rect 1409 6273 1443 6307
rect 5549 6273 5583 6307
rect 6929 6273 6963 6307
rect 7113 6273 7147 6307
rect 7389 6273 7423 6307
rect 7665 6273 7699 6307
rect 2697 6137 2731 6171
rect 7573 6137 7607 6171
rect 2053 6069 2087 6103
rect 4537 6069 4571 6103
rect 4905 6069 4939 6103
rect 5089 6069 5123 6103
rect 7021 6069 7055 6103
rect 7757 6069 7791 6103
rect 2145 5865 2179 5899
rect 4629 5865 4663 5899
rect 6653 5865 6687 5899
rect 7297 5865 7331 5899
rect 7481 5865 7515 5899
rect 4353 5797 4387 5831
rect 1501 5729 1535 5763
rect 7665 5729 7699 5763
rect 7941 5729 7975 5763
rect 1777 5661 1811 5695
rect 2237 5661 2271 5695
rect 2329 5661 2363 5695
rect 3985 5661 4019 5695
rect 6929 5661 6963 5695
rect 7389 5661 7423 5695
rect 7757 5661 7791 5695
rect 7849 5661 7883 5695
rect 4169 5593 4203 5627
rect 4813 5593 4847 5627
rect 7113 5593 7147 5627
rect 2421 5525 2455 5559
rect 4445 5525 4479 5559
rect 4613 5525 4647 5559
rect 7021 5525 7055 5559
rect 4077 5321 4111 5355
rect 4261 5321 4295 5355
rect 7021 5321 7055 5355
rect 7205 5321 7239 5355
rect 1777 5253 1811 5287
rect 4629 5253 4663 5287
rect 6469 5253 6503 5287
rect 3709 5185 3743 5219
rect 6377 5185 6411 5219
rect 7202 5185 7236 5219
rect 8033 5185 8067 5219
rect 1501 5117 1535 5151
rect 4353 5117 4387 5151
rect 6101 5117 6135 5151
rect 7665 5117 7699 5151
rect 3249 5049 3283 5083
rect 7849 5049 7883 5083
rect 4077 4981 4111 5015
rect 7573 4981 7607 5015
rect 2053 4777 2087 4811
rect 2237 4777 2271 4811
rect 3157 4777 3191 4811
rect 3893 4777 3927 4811
rect 5549 4777 5583 4811
rect 7757 4777 7791 4811
rect 2605 4709 2639 4743
rect 7205 4641 7239 4675
rect 7573 4641 7607 4675
rect 3341 4573 3375 4607
rect 3525 4573 3559 4607
rect 4261 4573 4295 4607
rect 5641 4573 5675 4607
rect 6929 4573 6963 4607
rect 7481 4573 7515 4607
rect 2237 4505 2271 4539
rect 4077 4505 4111 4539
rect 7113 4505 7147 4539
rect 6377 4437 6411 4471
rect 2697 4097 2731 4131
rect 3157 4097 3191 4131
rect 3801 4097 3835 4131
rect 3985 4097 4019 4131
rect 4445 4097 4479 4131
rect 6377 4097 6411 4131
rect 7021 4097 7055 4131
rect 7114 4097 7148 4131
rect 2053 4029 2087 4063
rect 3065 4029 3099 4063
rect 4721 4029 4755 4063
rect 6193 4029 6227 4063
rect 2881 3893 2915 3927
rect 3893 3893 3927 3927
rect 6469 3893 6503 3927
rect 7205 3893 7239 3927
rect 1409 3689 1443 3723
rect 3433 3689 3467 3723
rect 5917 3689 5951 3723
rect 6285 3689 6319 3723
rect 6745 3689 6779 3723
rect 7665 3689 7699 3723
rect 5089 3621 5123 3655
rect 7849 3621 7883 3655
rect 2881 3553 2915 3587
rect 3157 3553 3191 3587
rect 6101 3553 6135 3587
rect 6561 3553 6595 3587
rect 3801 3485 3835 3519
rect 5641 3485 5675 3519
rect 5733 3485 5767 3519
rect 6377 3485 6411 3519
rect 7021 3485 7055 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 8033 3485 8067 3519
rect 3249 3417 3283 3451
rect 6929 3417 6963 3451
rect 7113 3417 7147 3451
rect 3449 3349 3483 3383
rect 3617 3349 3651 3383
rect 7481 3349 7515 3383
rect 1501 3145 1535 3179
rect 2237 3145 2271 3179
rect 3985 3145 4019 3179
rect 6193 3145 6227 3179
rect 7389 3145 7423 3179
rect 4169 3077 4203 3111
rect 4721 3077 4755 3111
rect 6469 3077 6503 3111
rect 7297 3077 7331 3111
rect 1685 3009 1719 3043
rect 2145 3009 2179 3043
rect 4353 3009 4387 3043
rect 4445 3009 4479 3043
rect 6377 3009 6411 3043
rect 6929 3009 6963 3043
rect 7022 3009 7056 3043
rect 7603 3009 7637 3043
rect 7757 3009 7791 3043
rect 8033 3009 8067 3043
rect 7849 2805 7883 2839
rect 7481 2533 7515 2567
rect 7113 2397 7147 2431
rect 7267 2397 7301 2431
<< metal1 >>
rect 1104 9274 8372 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 8372 9274
rect 1104 9200 8372 9222
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4120 9132 5120 9160
rect 4120 9120 4126 9132
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 3881 9095 3939 9101
rect 3881 9092 3893 9095
rect 3844 9064 3893 9092
rect 3844 9052 3850 9064
rect 3881 9061 3893 9064
rect 3927 9092 3939 9095
rect 3927 9064 4752 9092
rect 3927 9061 3939 9064
rect 3881 9055 3939 9061
rect 4724 8965 4752 9064
rect 4616 8959 4674 8965
rect 4616 8956 4628 8959
rect 4595 8928 4628 8956
rect 4616 8925 4628 8928
rect 4662 8925 4674 8959
rect 4616 8919 4674 8925
rect 4709 8959 4767 8965
rect 4709 8925 4721 8959
rect 4755 8925 4767 8959
rect 4709 8919 4767 8925
rect 3142 8848 3148 8900
rect 3200 8888 3206 8900
rect 3329 8891 3387 8897
rect 3329 8888 3341 8891
rect 3200 8860 3341 8888
rect 3200 8848 3206 8860
rect 3329 8857 3341 8860
rect 3375 8857 3387 8891
rect 3329 8851 3387 8857
rect 4249 8891 4307 8897
rect 4249 8857 4261 8891
rect 4295 8888 4307 8891
rect 4632 8888 4660 8919
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4856 8928 4997 8956
rect 4856 8916 4862 8928
rect 4985 8925 4997 8928
rect 5031 8925 5043 8959
rect 5092 8956 5120 9132
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 5092 8928 5273 8956
rect 4985 8919 5043 8925
rect 5261 8925 5273 8928
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 4295 8860 5120 8888
rect 4295 8857 4307 8860
rect 4249 8851 4307 8857
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 4062 8820 4068 8832
rect 3835 8792 4068 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4341 8823 4399 8829
rect 4341 8789 4353 8823
rect 4387 8820 4399 8823
rect 4706 8820 4712 8832
rect 4387 8792 4712 8820
rect 4387 8789 4399 8792
rect 4341 8783 4399 8789
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 4798 8780 4804 8832
rect 4856 8780 4862 8832
rect 5092 8829 5120 8860
rect 5077 8823 5135 8829
rect 5077 8789 5089 8823
rect 5123 8789 5135 8823
rect 5077 8783 5135 8789
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 6733 8823 6791 8829
rect 6733 8820 6745 8823
rect 6696 8792 6745 8820
rect 6696 8780 6702 8792
rect 6733 8789 6745 8792
rect 6779 8789 6791 8823
rect 6733 8783 6791 8789
rect 1104 8730 8372 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 8372 8730
rect 1104 8656 8372 8678
rect 4341 8551 4399 8557
rect 4341 8517 4353 8551
rect 4387 8548 4399 8551
rect 4614 8548 4620 8560
rect 4387 8520 4620 8548
rect 4387 8517 4399 8520
rect 4341 8511 4399 8517
rect 4614 8508 4620 8520
rect 4672 8508 4678 8560
rect 5718 8508 5724 8560
rect 5776 8508 5782 8560
rect 7193 8551 7251 8557
rect 7193 8548 7205 8551
rect 6656 8520 7205 8548
rect 6656 8492 6684 8520
rect 7193 8517 7205 8520
rect 7239 8517 7251 8551
rect 7193 8511 7251 8517
rect 6638 8440 6644 8492
rect 6696 8440 6702 8492
rect 6734 8483 6792 8489
rect 6734 8449 6746 8483
rect 6780 8449 6792 8483
rect 6734 8443 6792 8449
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 4433 8415 4491 8421
rect 4433 8412 4445 8415
rect 3200 8384 4445 8412
rect 3200 8372 3206 8384
rect 4433 8381 4445 8384
rect 4479 8381 4491 8415
rect 4433 8375 4491 8381
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 4798 8412 4804 8424
rect 4755 8384 4804 8412
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 4798 8372 4804 8384
rect 4856 8372 4862 8424
rect 6748 8412 6776 8443
rect 6822 8440 6828 8492
rect 6880 8480 6886 8492
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6880 8452 7113 8480
rect 6880 8440 6886 8452
rect 7101 8449 7113 8452
rect 7147 8449 7159 8483
rect 7101 8443 7159 8449
rect 7377 8483 7435 8489
rect 7377 8449 7389 8483
rect 7423 8480 7435 8483
rect 7466 8480 7472 8492
rect 7423 8452 7472 8480
rect 7423 8449 7435 8452
rect 7377 8443 7435 8449
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 6196 8384 6776 8412
rect 6196 8288 6224 8384
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7009 8347 7067 8353
rect 7009 8344 7021 8347
rect 6972 8316 7021 8344
rect 6972 8304 6978 8316
rect 7009 8313 7021 8316
rect 7055 8313 7067 8347
rect 7009 8307 7067 8313
rect 3053 8279 3111 8285
rect 3053 8245 3065 8279
rect 3099 8276 3111 8279
rect 3142 8276 3148 8288
rect 3099 8248 3148 8276
rect 3099 8245 3111 8248
rect 3053 8239 3111 8245
rect 3142 8236 3148 8248
rect 3200 8236 3206 8288
rect 3878 8236 3884 8288
rect 3936 8276 3942 8288
rect 6086 8276 6092 8288
rect 3936 8248 6092 8276
rect 3936 8236 3942 8248
rect 6086 8236 6092 8248
rect 6144 8236 6150 8288
rect 6178 8236 6184 8288
rect 6236 8236 6242 8288
rect 7374 8236 7380 8288
rect 7432 8236 7438 8288
rect 1104 8186 8372 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 8372 8186
rect 1104 8112 8372 8134
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 3108 8044 3433 8072
rect 3108 8032 3114 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3421 8035 3479 8041
rect 3786 8032 3792 8084
rect 3844 8072 3850 8084
rect 4709 8075 4767 8081
rect 4709 8072 4721 8075
rect 3844 8044 4721 8072
rect 3844 8032 3850 8044
rect 4709 8041 4721 8044
rect 4755 8041 4767 8075
rect 4709 8035 4767 8041
rect 5718 8032 5724 8084
rect 5776 8032 5782 8084
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 6822 8072 6828 8084
rect 6052 8044 6828 8072
rect 6052 8032 6058 8044
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 3878 7964 3884 8016
rect 3936 7964 3942 8016
rect 4246 7964 4252 8016
rect 4304 8004 4310 8016
rect 4890 8004 4896 8016
rect 4304 7976 4896 8004
rect 4304 7964 4310 7976
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 7469 8007 7527 8013
rect 7469 8004 7481 8007
rect 6886 7976 7481 8004
rect 4706 7936 4712 7948
rect 4172 7908 4712 7936
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 2222 7760 2228 7812
rect 2280 7760 2286 7812
rect 2869 7803 2927 7809
rect 2869 7769 2881 7803
rect 2915 7800 2927 7803
rect 3605 7803 3663 7809
rect 2915 7772 3280 7800
rect 2915 7769 2927 7772
rect 2869 7763 2927 7769
rect 1397 7735 1455 7741
rect 1397 7701 1409 7735
rect 1443 7732 1455 7735
rect 2774 7732 2780 7744
rect 1443 7704 2780 7732
rect 1443 7701 1455 7704
rect 1397 7695 1455 7701
rect 2774 7692 2780 7704
rect 2832 7692 2838 7744
rect 3252 7741 3280 7772
rect 3605 7769 3617 7803
rect 3651 7769 3663 7803
rect 4172 7800 4200 7908
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 5994 7936 6000 7948
rect 5184 7908 6000 7936
rect 4341 7849 4399 7855
rect 4341 7815 4353 7849
rect 4387 7846 4399 7849
rect 4387 7818 4476 7846
rect 4522 7828 4528 7880
rect 4580 7828 4586 7880
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 5074 7868 5080 7880
rect 5031 7840 5080 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 5074 7828 5080 7840
rect 5132 7828 5138 7880
rect 5184 7877 5212 7908
rect 5994 7896 6000 7908
rect 6052 7896 6058 7948
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6641 7939 6699 7945
rect 6144 7908 6316 7936
rect 6144 7896 6150 7908
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5776 7840 5825 7868
rect 5776 7828 5782 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 5905 7871 5963 7877
rect 5905 7837 5917 7871
rect 5951 7868 5963 7871
rect 6178 7868 6184 7880
rect 5951 7840 6184 7868
rect 5951 7837 5963 7840
rect 5905 7831 5963 7837
rect 4387 7815 4399 7818
rect 4341 7809 4399 7815
rect 4249 7803 4307 7809
rect 4249 7800 4261 7803
rect 4172 7772 4261 7800
rect 3605 7763 3663 7769
rect 4249 7769 4261 7772
rect 4295 7769 4307 7803
rect 4249 7763 4307 7769
rect 3418 7741 3424 7744
rect 3237 7735 3295 7741
rect 3237 7701 3249 7735
rect 3283 7701 3295 7735
rect 3237 7695 3295 7701
rect 3405 7735 3424 7741
rect 3405 7701 3417 7735
rect 3405 7695 3424 7701
rect 3418 7692 3424 7695
rect 3476 7692 3482 7744
rect 3620 7732 3648 7763
rect 4448 7744 4476 7818
rect 4540 7800 4568 7828
rect 4677 7803 4735 7809
rect 4677 7800 4689 7803
rect 4540 7772 4689 7800
rect 4677 7769 4689 7772
rect 4723 7769 4735 7803
rect 4677 7763 4735 7769
rect 4893 7803 4951 7809
rect 4893 7769 4905 7803
rect 4939 7800 4951 7803
rect 5920 7800 5948 7831
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6288 7868 6316 7908
rect 6641 7905 6653 7939
rect 6687 7936 6699 7939
rect 6886 7936 6914 7976
rect 7469 7973 7481 7976
rect 7515 7973 7527 8007
rect 7469 7967 7527 7973
rect 6687 7908 6914 7936
rect 7101 7939 7159 7945
rect 6687 7905 6699 7908
rect 6641 7899 6699 7905
rect 7101 7905 7113 7939
rect 7147 7936 7159 7939
rect 7374 7936 7380 7948
rect 7147 7908 7380 7936
rect 7147 7905 7159 7908
rect 7101 7899 7159 7905
rect 7374 7896 7380 7908
rect 7432 7896 7438 7948
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6288 7840 6745 7868
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 6733 7831 6791 7837
rect 7024 7840 7205 7868
rect 4939 7772 5948 7800
rect 4939 7769 4951 7772
rect 4893 7763 4951 7769
rect 7024 7744 7052 7840
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 7098 7760 7104 7812
rect 7156 7800 7162 7812
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 7156 7772 7297 7800
rect 7156 7760 7162 7772
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7285 7763 7343 7769
rect 4154 7732 4160 7744
rect 3620 7704 4160 7732
rect 4154 7692 4160 7704
rect 4212 7692 4218 7744
rect 4430 7692 4436 7744
rect 4488 7692 4494 7744
rect 4522 7692 4528 7744
rect 4580 7692 4586 7744
rect 4798 7692 4804 7744
rect 4856 7732 4862 7744
rect 5077 7735 5135 7741
rect 5077 7732 5089 7735
rect 4856 7704 5089 7732
rect 4856 7692 4862 7704
rect 5077 7701 5089 7704
rect 5123 7701 5135 7735
rect 5077 7695 5135 7701
rect 6457 7735 6515 7741
rect 6457 7701 6469 7735
rect 6503 7732 6515 7735
rect 6730 7732 6736 7744
rect 6503 7704 6736 7732
rect 6503 7701 6515 7704
rect 6457 7695 6515 7701
rect 6730 7692 6736 7704
rect 6788 7692 6794 7744
rect 6914 7692 6920 7744
rect 6972 7692 6978 7744
rect 7006 7692 7012 7744
rect 7064 7692 7070 7744
rect 1104 7642 8372 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 8372 7642
rect 1104 7568 8372 7590
rect 2222 7488 2228 7540
rect 2280 7488 2286 7540
rect 3050 7488 3056 7540
rect 3108 7488 3114 7540
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 5258 7528 5264 7540
rect 4540 7500 5264 7528
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 2869 7463 2927 7469
rect 2869 7460 2881 7463
rect 2832 7432 2881 7460
rect 2832 7420 2838 7432
rect 2869 7429 2881 7432
rect 2915 7429 2927 7463
rect 2869 7423 2927 7429
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2406 7392 2412 7404
rect 2363 7364 2412 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2406 7352 2412 7364
rect 2464 7352 2470 7404
rect 2682 7352 2688 7404
rect 2740 7352 2746 7404
rect 2884 7392 2912 7423
rect 3418 7420 3424 7472
rect 3476 7460 3482 7472
rect 3881 7463 3939 7469
rect 3881 7460 3893 7463
rect 3476 7432 3893 7460
rect 3476 7420 3482 7432
rect 3881 7429 3893 7432
rect 3927 7460 3939 7463
rect 4540 7460 4568 7500
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 6825 7531 6883 7537
rect 6825 7497 6837 7531
rect 6871 7528 6883 7531
rect 7006 7528 7012 7540
rect 6871 7500 7012 7528
rect 6871 7497 6883 7500
rect 6825 7491 6883 7497
rect 7006 7488 7012 7500
rect 7064 7488 7070 7540
rect 7285 7531 7343 7537
rect 7285 7497 7297 7531
rect 7331 7528 7343 7531
rect 7466 7528 7472 7540
rect 7331 7500 7472 7528
rect 7331 7497 7343 7500
rect 7285 7491 7343 7497
rect 7466 7488 7472 7500
rect 7524 7488 7530 7540
rect 3927 7432 4568 7460
rect 4709 7463 4767 7469
rect 3927 7429 3939 7432
rect 3881 7423 3939 7429
rect 4709 7429 4721 7463
rect 4755 7460 4767 7463
rect 4890 7460 4896 7472
rect 4755 7432 4896 7460
rect 4755 7429 4767 7432
rect 4709 7423 4767 7429
rect 4890 7420 4896 7432
rect 4948 7420 4954 7472
rect 3786 7392 3792 7404
rect 2884 7364 3792 7392
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 4246 7401 4252 7404
rect 3973 7395 4031 7401
rect 3973 7361 3985 7395
rect 4019 7392 4031 7395
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 4019 7364 4077 7392
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 4219 7395 4252 7401
rect 4219 7361 4231 7395
rect 4219 7355 4252 7361
rect 2700 7324 2728 7352
rect 3988 7324 4016 7355
rect 4246 7352 4252 7355
rect 4304 7352 4310 7404
rect 4522 7352 4528 7404
rect 4580 7392 4586 7404
rect 5077 7395 5135 7401
rect 5077 7392 5089 7395
rect 4580 7364 5089 7392
rect 4580 7352 4586 7364
rect 5077 7361 5089 7364
rect 5123 7392 5135 7395
rect 5258 7392 5264 7404
rect 5123 7364 5264 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5258 7352 5264 7364
rect 5316 7352 5322 7404
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 7039 7395 7097 7401
rect 7039 7392 7051 7395
rect 6328 7364 7051 7392
rect 6328 7352 6334 7364
rect 7024 7361 7051 7364
rect 7085 7392 7097 7395
rect 7193 7395 7251 7401
rect 7085 7364 7157 7392
rect 7085 7361 7097 7364
rect 7024 7355 7097 7361
rect 7193 7361 7205 7395
rect 7239 7392 7251 7395
rect 7239 7364 7880 7392
rect 7239 7361 7251 7364
rect 7193 7355 7251 7361
rect 4338 7324 4344 7336
rect 2700 7296 4344 7324
rect 4338 7284 4344 7296
rect 4396 7284 4402 7336
rect 4706 7324 4712 7336
rect 4540 7296 4712 7324
rect 4540 7265 4568 7296
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 7024 7324 7052 7355
rect 7745 7327 7803 7333
rect 7745 7324 7757 7327
rect 7024 7296 7757 7324
rect 7745 7293 7757 7296
rect 7791 7293 7803 7327
rect 7745 7287 7803 7293
rect 4525 7259 4583 7265
rect 4525 7225 4537 7259
rect 4571 7225 4583 7259
rect 4890 7256 4896 7268
rect 4525 7219 4583 7225
rect 4632 7228 4896 7256
rect 4154 7148 4160 7200
rect 4212 7188 4218 7200
rect 4632 7188 4660 7228
rect 4890 7216 4896 7228
rect 4948 7216 4954 7268
rect 7852 7265 7880 7364
rect 8018 7352 8024 7404
rect 8076 7352 8082 7404
rect 7469 7259 7527 7265
rect 7469 7225 7481 7259
rect 7515 7256 7527 7259
rect 7837 7259 7895 7265
rect 7837 7256 7849 7259
rect 7515 7228 7849 7256
rect 7515 7225 7527 7228
rect 7469 7219 7527 7225
rect 7837 7225 7849 7228
rect 7883 7225 7895 7259
rect 7837 7219 7895 7225
rect 4212 7160 4660 7188
rect 4709 7191 4767 7197
rect 4212 7148 4218 7160
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 4798 7188 4804 7200
rect 4755 7160 4804 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 1104 7098 8372 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 8372 7098
rect 1104 7024 8372 7046
rect 4249 6987 4307 6993
rect 4249 6953 4261 6987
rect 4295 6984 4307 6987
rect 4798 6984 4804 6996
rect 4295 6956 4804 6984
rect 4295 6953 4307 6956
rect 4249 6947 4307 6953
rect 4798 6944 4804 6956
rect 4856 6944 4862 6996
rect 4433 6919 4491 6925
rect 4433 6885 4445 6919
rect 4479 6916 4491 6919
rect 4479 6888 4660 6916
rect 4479 6885 4491 6888
rect 4433 6879 4491 6885
rect 3142 6808 3148 6860
rect 3200 6848 3206 6860
rect 4525 6851 4583 6857
rect 4525 6848 4537 6851
rect 3200 6820 4537 6848
rect 3200 6808 3206 6820
rect 4525 6817 4537 6820
rect 4571 6817 4583 6851
rect 4632 6848 4660 6888
rect 4801 6851 4859 6857
rect 4801 6848 4813 6851
rect 4632 6820 4813 6848
rect 4525 6811 4583 6817
rect 4801 6817 4813 6820
rect 4847 6817 4859 6851
rect 4801 6811 4859 6817
rect 4890 6808 4896 6860
rect 4948 6848 4954 6860
rect 6086 6848 6092 6860
rect 4948 6820 6092 6848
rect 4948 6808 4954 6820
rect 6086 6808 6092 6820
rect 6144 6848 6150 6860
rect 6144 6820 6914 6848
rect 6144 6808 6150 6820
rect 3326 6740 3332 6792
rect 3384 6740 3390 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3421 6743 3479 6749
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6749 3939 6783
rect 3881 6743 3939 6749
rect 2130 6672 2136 6724
rect 2188 6672 2194 6724
rect 2866 6672 2872 6724
rect 2924 6672 2930 6724
rect 1397 6647 1455 6653
rect 1397 6613 1409 6647
rect 1443 6644 1455 6647
rect 2682 6644 2688 6656
rect 1443 6616 2688 6644
rect 1443 6613 1455 6616
rect 1397 6607 1455 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 3436 6644 3464 6743
rect 3605 6715 3663 6721
rect 3605 6681 3617 6715
rect 3651 6712 3663 6715
rect 3896 6712 3924 6743
rect 6638 6740 6644 6792
rect 6696 6740 6702 6792
rect 6730 6740 6736 6792
rect 6788 6740 6794 6792
rect 4706 6712 4712 6724
rect 3651 6684 4712 6712
rect 3651 6681 3663 6684
rect 3605 6675 3663 6681
rect 4706 6672 4712 6684
rect 4764 6672 4770 6724
rect 5534 6672 5540 6724
rect 5592 6672 5598 6724
rect 4154 6644 4160 6656
rect 3436 6616 4160 6644
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 4890 6644 4896 6656
rect 4304 6616 4896 6644
rect 4304 6604 4310 6616
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 6270 6604 6276 6656
rect 6328 6604 6334 6656
rect 6886 6644 6914 6820
rect 7466 6740 7472 6792
rect 7524 6740 7530 6792
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 6886 6616 7389 6644
rect 7377 6613 7389 6616
rect 7423 6613 7435 6647
rect 7377 6607 7435 6613
rect 1104 6554 8372 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 8372 6554
rect 1104 6480 8372 6502
rect 2777 6443 2835 6449
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 2866 6440 2872 6452
rect 2823 6412 2872 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 2866 6400 2872 6412
rect 2924 6400 2930 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5629 6443 5687 6449
rect 5629 6440 5641 6443
rect 5592 6412 5641 6440
rect 5592 6400 5598 6412
rect 5629 6409 5641 6412
rect 5675 6409 5687 6443
rect 5629 6403 5687 6409
rect 2317 6375 2375 6381
rect 2317 6341 2329 6375
rect 2363 6372 2375 6375
rect 2682 6372 2688 6384
rect 2363 6344 2688 6372
rect 2363 6341 2375 6344
rect 2317 6335 2375 6341
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 3050 6332 3056 6384
rect 3108 6332 3114 6384
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 5061 6375 5119 6381
rect 5061 6372 5073 6375
rect 4212 6344 5073 6372
rect 4212 6332 4218 6344
rect 5061 6341 5073 6344
rect 5107 6372 5119 6375
rect 5166 6372 5172 6384
rect 5107 6344 5172 6372
rect 5107 6341 5119 6344
rect 5061 6335 5119 6341
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 5261 6375 5319 6381
rect 5261 6341 5273 6375
rect 5307 6372 5319 6375
rect 5350 6372 5356 6384
rect 5307 6344 5356 6372
rect 5307 6341 5319 6344
rect 5261 6335 5319 6341
rect 5350 6332 5356 6344
rect 5408 6332 5414 6384
rect 842 6264 848 6316
rect 900 6304 906 6316
rect 1397 6307 1455 6313
rect 1397 6304 1409 6307
rect 900 6276 1409 6304
rect 900 6264 906 6276
rect 1397 6273 1409 6276
rect 1443 6273 1455 6307
rect 1397 6267 1455 6273
rect 2406 6264 2412 6316
rect 2464 6304 2470 6316
rect 5534 6304 5540 6316
rect 2464 6276 5540 6304
rect 2464 6264 2470 6276
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 6917 6307 6975 6313
rect 6917 6273 6929 6307
rect 6963 6304 6975 6307
rect 7006 6304 7012 6316
rect 6963 6276 7012 6304
rect 6963 6273 6975 6276
rect 6917 6267 6975 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7098 6264 7104 6316
rect 7156 6264 7162 6316
rect 7374 6264 7380 6316
rect 7432 6264 7438 6316
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7576 6276 7665 6304
rect 2685 6171 2743 6177
rect 2685 6137 2697 6171
rect 2731 6137 2743 6171
rect 2685 6131 2743 6137
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 2041 6103 2099 6109
rect 2041 6100 2053 6103
rect 1820 6072 2053 6100
rect 1820 6060 1826 6072
rect 2041 6069 2053 6072
rect 2087 6069 2099 6103
rect 2041 6063 2099 6069
rect 2222 6060 2228 6112
rect 2280 6100 2286 6112
rect 2700 6100 2728 6131
rect 3326 6128 3332 6180
rect 3384 6168 3390 6180
rect 6270 6168 6276 6180
rect 3384 6140 6276 6168
rect 3384 6128 3390 6140
rect 3970 6100 3976 6112
rect 2280 6072 3976 6100
rect 2280 6060 2286 6072
rect 3970 6060 3976 6072
rect 4028 6100 4034 6112
rect 4246 6100 4252 6112
rect 4028 6072 4252 6100
rect 4028 6060 4034 6072
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 4525 6103 4583 6109
rect 4525 6069 4537 6103
rect 4571 6100 4583 6103
rect 4614 6100 4620 6112
rect 4571 6072 4620 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 4890 6060 4896 6112
rect 4948 6060 4954 6112
rect 5092 6109 5120 6140
rect 6270 6128 6276 6140
rect 6328 6128 6334 6180
rect 7576 6177 7604 6276
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 7653 6267 7711 6273
rect 7561 6171 7619 6177
rect 7561 6137 7573 6171
rect 7607 6137 7619 6171
rect 7561 6131 7619 6137
rect 5077 6103 5135 6109
rect 5077 6069 5089 6103
rect 5123 6069 5135 6103
rect 5077 6063 5135 6069
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7009 6103 7067 6109
rect 7009 6100 7021 6103
rect 6972 6072 7021 6100
rect 6972 6060 6978 6072
rect 7009 6069 7021 6072
rect 7055 6069 7067 6103
rect 7009 6063 7067 6069
rect 7282 6060 7288 6112
rect 7340 6100 7346 6112
rect 7745 6103 7803 6109
rect 7745 6100 7757 6103
rect 7340 6072 7757 6100
rect 7340 6060 7346 6072
rect 7745 6069 7757 6072
rect 7791 6069 7803 6103
rect 7745 6063 7803 6069
rect 1104 6010 8372 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 8372 6010
rect 1104 5936 8372 5958
rect 2130 5856 2136 5908
rect 2188 5856 2194 5908
rect 4617 5899 4675 5905
rect 4617 5865 4629 5899
rect 4663 5896 4675 5899
rect 5350 5896 5356 5908
rect 4663 5868 5356 5896
rect 4663 5865 4675 5868
rect 4617 5859 4675 5865
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 6638 5856 6644 5908
rect 6696 5856 6702 5908
rect 7282 5856 7288 5908
rect 7340 5856 7346 5908
rect 7466 5856 7472 5908
rect 7524 5856 7530 5908
rect 4341 5831 4399 5837
rect 4341 5797 4353 5831
rect 4387 5828 4399 5831
rect 4798 5828 4804 5840
rect 4387 5800 4804 5828
rect 4387 5797 4399 5800
rect 4341 5791 4399 5797
rect 4798 5788 4804 5800
rect 4856 5788 4862 5840
rect 6730 5788 6736 5840
rect 6788 5828 6794 5840
rect 6788 5800 7972 5828
rect 6788 5788 6794 5800
rect 1489 5763 1547 5769
rect 1489 5729 1501 5763
rect 1535 5760 1547 5763
rect 1535 5732 2268 5760
rect 1535 5729 1547 5732
rect 1489 5723 1547 5729
rect 1762 5652 1768 5704
rect 1820 5652 1826 5704
rect 2240 5701 2268 5732
rect 4154 5720 4160 5772
rect 4212 5760 4218 5772
rect 4890 5760 4896 5772
rect 4212 5732 4896 5760
rect 4212 5720 4218 5732
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 7944 5769 7972 5800
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 6932 5732 7665 5760
rect 6932 5704 6960 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5692 2283 5695
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2271 5664 2329 5692
rect 2271 5661 2283 5664
rect 2225 5655 2283 5661
rect 2317 5661 2329 5664
rect 2363 5692 2375 5695
rect 2406 5692 2412 5704
rect 2363 5664 2412 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4062 5692 4068 5704
rect 4019 5664 4068 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 7742 5652 7748 5704
rect 7800 5652 7806 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 3326 5584 3332 5636
rect 3384 5624 3390 5636
rect 4157 5627 4215 5633
rect 4157 5624 4169 5627
rect 3384 5596 4169 5624
rect 3384 5584 3390 5596
rect 4157 5593 4169 5596
rect 4203 5593 4215 5627
rect 4157 5587 4215 5593
rect 4246 5584 4252 5636
rect 4304 5624 4310 5636
rect 4801 5627 4859 5633
rect 4801 5624 4813 5627
rect 4304 5596 4813 5624
rect 4304 5584 4310 5596
rect 4801 5593 4813 5596
rect 4847 5624 4859 5627
rect 5258 5624 5264 5636
rect 4847 5596 5264 5624
rect 4847 5593 4859 5596
rect 4801 5587 4859 5593
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 7024 5624 7052 5652
rect 6932 5596 7052 5624
rect 7101 5627 7159 5633
rect 6932 5568 6960 5596
rect 7101 5593 7113 5627
rect 7147 5624 7159 5627
rect 7650 5624 7656 5636
rect 7147 5596 7656 5624
rect 7147 5593 7159 5596
rect 7101 5587 7159 5593
rect 7650 5584 7656 5596
rect 7708 5624 7714 5636
rect 7852 5624 7880 5655
rect 7708 5596 7880 5624
rect 7708 5584 7714 5596
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 2774 5556 2780 5568
rect 2455 5528 2780 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 2774 5516 2780 5528
rect 2832 5516 2838 5568
rect 3786 5516 3792 5568
rect 3844 5556 3850 5568
rect 4433 5559 4491 5565
rect 4433 5556 4445 5559
rect 3844 5528 4445 5556
rect 3844 5516 3850 5528
rect 4433 5525 4445 5528
rect 4479 5525 4491 5559
rect 4433 5519 4491 5525
rect 4601 5559 4659 5565
rect 4601 5525 4613 5559
rect 4647 5556 4659 5559
rect 4706 5556 4712 5568
rect 4647 5528 4712 5556
rect 4647 5525 4659 5528
rect 4601 5519 4659 5525
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 6914 5516 6920 5568
rect 6972 5516 6978 5568
rect 7006 5516 7012 5568
rect 7064 5516 7070 5568
rect 1104 5466 8372 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 8372 5466
rect 1104 5392 8372 5414
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 4065 5355 4123 5361
rect 4065 5352 4077 5355
rect 4028 5324 4077 5352
rect 4028 5312 4034 5324
rect 4065 5321 4077 5324
rect 4111 5321 4123 5355
rect 4065 5315 4123 5321
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4295 5324 4660 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 2038 5284 2044 5296
rect 1811 5256 2044 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 2038 5244 2044 5256
rect 2096 5244 2102 5296
rect 2774 5244 2780 5296
rect 2832 5244 2838 5296
rect 4632 5293 4660 5324
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 5316 5324 6408 5352
rect 5316 5312 5322 5324
rect 4617 5287 4675 5293
rect 4617 5253 4629 5287
rect 4663 5253 4675 5287
rect 4617 5247 4675 5253
rect 5626 5244 5632 5296
rect 5684 5244 5690 5296
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5216 3755 5219
rect 4154 5216 4160 5228
rect 3743 5188 4160 5216
rect 3743 5185 3755 5188
rect 3697 5179 3755 5185
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 6380 5225 6408 5324
rect 7006 5312 7012 5364
rect 7064 5312 7070 5364
rect 7193 5355 7251 5361
rect 7193 5321 7205 5355
rect 7239 5352 7251 5355
rect 7282 5352 7288 5364
rect 7239 5324 7288 5352
rect 7239 5321 7251 5324
rect 7193 5315 7251 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 6457 5287 6515 5293
rect 6457 5253 6469 5287
rect 6503 5284 6515 5287
rect 6914 5284 6920 5296
rect 6503 5256 6920 5284
rect 6503 5253 6515 5256
rect 6457 5247 6515 5253
rect 6914 5244 6920 5256
rect 6972 5244 6978 5296
rect 6365 5219 6423 5225
rect 6365 5185 6377 5219
rect 6411 5185 6423 5219
rect 7190 5219 7248 5225
rect 7190 5216 7202 5219
rect 6365 5179 6423 5185
rect 6886 5188 7202 5216
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 1535 5120 4353 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 3237 5083 3295 5089
rect 3237 5049 3249 5083
rect 3283 5080 3295 5083
rect 3326 5080 3332 5092
rect 3283 5052 3332 5080
rect 3283 5049 3295 5052
rect 3237 5043 3295 5049
rect 3326 5040 3332 5052
rect 3384 5080 3390 5092
rect 4246 5080 4252 5092
rect 3384 5052 4252 5080
rect 3384 5040 3390 5052
rect 4246 5040 4252 5052
rect 4304 5040 4310 5092
rect 3878 4972 3884 5024
rect 3936 5012 3942 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 3936 4984 4077 5012
rect 3936 4972 3942 4984
rect 4065 4981 4077 4984
rect 4111 4981 4123 5015
rect 4356 5012 4384 5111
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 6089 5151 6147 5157
rect 6089 5148 6101 5151
rect 5408 5120 6101 5148
rect 5408 5108 5414 5120
rect 6089 5117 6101 5120
rect 6135 5148 6147 5151
rect 6886 5148 6914 5188
rect 7190 5185 7202 5188
rect 7236 5216 7248 5219
rect 7374 5216 7380 5228
rect 7236 5188 7380 5216
rect 7236 5185 7248 5188
rect 7190 5179 7248 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 8018 5176 8024 5228
rect 8076 5176 8082 5228
rect 6135 5120 6914 5148
rect 6135 5117 6147 5120
rect 6089 5111 6147 5117
rect 7098 5108 7104 5160
rect 7156 5148 7162 5160
rect 7558 5148 7564 5160
rect 7156 5120 7564 5148
rect 7156 5108 7162 5120
rect 7558 5108 7564 5120
rect 7616 5148 7622 5160
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7616 5120 7665 5148
rect 7616 5108 7622 5120
rect 7653 5117 7665 5120
rect 7699 5148 7711 5151
rect 7699 5120 7880 5148
rect 7699 5117 7711 5120
rect 7653 5111 7711 5117
rect 7852 5089 7880 5120
rect 7837 5083 7895 5089
rect 7837 5049 7849 5083
rect 7883 5049 7895 5083
rect 7837 5043 7895 5049
rect 4706 5012 4712 5024
rect 4356 4984 4712 5012
rect 4065 4975 4123 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7466 5012 7472 5024
rect 6972 4984 7472 5012
rect 6972 4972 6978 4984
rect 7466 4972 7472 4984
rect 7524 5012 7530 5024
rect 7561 5015 7619 5021
rect 7561 5012 7573 5015
rect 7524 4984 7573 5012
rect 7524 4972 7530 4984
rect 7561 4981 7573 4984
rect 7607 4981 7619 5015
rect 7561 4975 7619 4981
rect 1104 4922 8372 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 8372 4922
rect 1104 4848 8372 4870
rect 2038 4768 2044 4820
rect 2096 4768 2102 4820
rect 2225 4811 2283 4817
rect 2225 4777 2237 4811
rect 2271 4808 2283 4811
rect 3145 4811 3203 4817
rect 3145 4808 3157 4811
rect 2271 4780 3157 4808
rect 2271 4777 2283 4780
rect 2225 4771 2283 4777
rect 3145 4777 3157 4780
rect 3191 4777 3203 4811
rect 3145 4771 3203 4777
rect 3878 4768 3884 4820
rect 3936 4768 3942 4820
rect 5537 4811 5595 4817
rect 5537 4777 5549 4811
rect 5583 4808 5595 4811
rect 5626 4808 5632 4820
rect 5583 4780 5632 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 5626 4768 5632 4780
rect 5684 4768 5690 4820
rect 7742 4768 7748 4820
rect 7800 4768 7806 4820
rect 2593 4743 2651 4749
rect 2593 4709 2605 4743
rect 2639 4740 2651 4743
rect 3786 4740 3792 4752
rect 2639 4712 3792 4740
rect 2639 4709 2651 4712
rect 2593 4703 2651 4709
rect 3786 4700 3792 4712
rect 3844 4700 3850 4752
rect 4062 4672 4068 4684
rect 3528 4644 4068 4672
rect 3326 4564 3332 4616
rect 3384 4564 3390 4616
rect 3528 4613 3556 4644
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 7193 4675 7251 4681
rect 7193 4641 7205 4675
rect 7239 4672 7251 4675
rect 7282 4672 7288 4684
rect 7239 4644 7288 4672
rect 7239 4641 7251 4644
rect 7193 4635 7251 4641
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 7558 4632 7564 4684
rect 7616 4632 7622 4684
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4573 3571 4607
rect 3513 4567 3571 4573
rect 4249 4607 4307 4613
rect 4249 4573 4261 4607
rect 4295 4604 4307 4607
rect 4798 4604 4804 4616
rect 4295 4576 4804 4604
rect 4295 4573 4307 4576
rect 4249 4567 4307 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 5534 4564 5540 4616
rect 5592 4604 5598 4616
rect 5629 4607 5687 4613
rect 5629 4604 5641 4607
rect 5592 4576 5641 4604
rect 5592 4564 5598 4576
rect 5629 4573 5641 4576
rect 5675 4604 5687 4607
rect 6178 4604 6184 4616
rect 5675 4576 6184 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 6178 4564 6184 4576
rect 6236 4564 6242 4616
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 7466 4564 7472 4616
rect 7524 4564 7530 4616
rect 2222 4496 2228 4548
rect 2280 4536 2286 4548
rect 3050 4536 3056 4548
rect 2280 4508 3056 4536
rect 2280 4496 2286 4508
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 4065 4539 4123 4545
rect 4065 4505 4077 4539
rect 4111 4536 4123 4539
rect 5350 4536 5356 4548
rect 4111 4508 5356 4536
rect 4111 4505 4123 4508
rect 4065 4499 4123 4505
rect 5350 4496 5356 4508
rect 5408 4536 5414 4548
rect 7101 4539 7159 4545
rect 7101 4536 7113 4539
rect 5408 4508 7113 4536
rect 5408 4496 5414 4508
rect 7101 4505 7113 4508
rect 7147 4505 7159 4539
rect 7101 4499 7159 4505
rect 6362 4428 6368 4480
rect 6420 4428 6426 4480
rect 1104 4378 8372 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 8372 4378
rect 1104 4304 8372 4326
rect 4706 4196 4712 4208
rect 4448 4168 4712 4196
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 3145 4131 3203 4137
rect 3145 4128 3157 4131
rect 2731 4100 3157 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 3145 4097 3157 4100
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3786 4088 3792 4140
rect 3844 4088 3850 4140
rect 3973 4131 4031 4137
rect 3973 4097 3985 4131
rect 4019 4128 4031 4131
rect 4062 4128 4068 4140
rect 4019 4100 4068 4128
rect 4019 4097 4031 4100
rect 3973 4091 4031 4097
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4448 4137 4476 4168
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 6270 4196 6276 4208
rect 5934 4168 6276 4196
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 4433 4131 4491 4137
rect 4433 4097 4445 4131
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 6362 4088 6368 4140
rect 6420 4088 6426 4140
rect 7006 4088 7012 4140
rect 7064 4088 7070 4140
rect 7102 4131 7160 4137
rect 7102 4097 7114 4131
rect 7148 4097 7160 4131
rect 7102 4091 7160 4097
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 2041 4063 2099 4069
rect 2041 4060 2053 4063
rect 1452 4032 2053 4060
rect 1452 4020 1458 4032
rect 2041 4029 2053 4032
rect 2087 4029 2099 4063
rect 2041 4023 2099 4029
rect 3050 4020 3056 4072
rect 3108 4020 3114 4072
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4060 4767 4063
rect 5902 4060 5908 4072
rect 4755 4032 5908 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6181 4063 6239 4069
rect 6181 4029 6193 4063
rect 6227 4060 6239 4063
rect 6914 4060 6920 4072
rect 6227 4032 6920 4060
rect 6227 4029 6239 4032
rect 6181 4023 6239 4029
rect 6914 4020 6920 4032
rect 6972 4060 6978 4072
rect 7116 4060 7144 4091
rect 6972 4032 7144 4060
rect 6972 4020 6978 4032
rect 2866 3884 2872 3936
rect 2924 3884 2930 3936
rect 3878 3884 3884 3936
rect 3936 3884 3942 3936
rect 5718 3884 5724 3936
rect 5776 3924 5782 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 5776 3896 6469 3924
rect 5776 3884 5782 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 6457 3887 6515 3893
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 7282 3924 7288 3936
rect 7239 3896 7288 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 1104 3834 8372 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 8372 3834
rect 1104 3760 8372 3782
rect 1394 3680 1400 3732
rect 1452 3680 1458 3732
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3720 3479 3723
rect 3878 3720 3884 3732
rect 3467 3692 3884 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 3878 3680 3884 3692
rect 3936 3720 3942 3732
rect 3936 3692 5672 3720
rect 3936 3680 3942 3692
rect 5077 3655 5135 3661
rect 5077 3652 5089 3655
rect 4724 3624 5089 3652
rect 4724 3596 4752 3624
rect 5077 3621 5089 3624
rect 5123 3621 5135 3655
rect 5077 3615 5135 3621
rect 2866 3544 2872 3596
rect 2924 3544 2930 3596
rect 3145 3587 3203 3593
rect 3145 3553 3157 3587
rect 3191 3584 3203 3587
rect 4430 3584 4436 3596
rect 3191 3556 4436 3584
rect 3191 3553 3203 3556
rect 3145 3547 3203 3553
rect 4430 3544 4436 3556
rect 4488 3584 4494 3596
rect 4706 3584 4712 3596
rect 4488 3556 4712 3584
rect 4488 3544 4494 3556
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 4614 3516 4620 3528
rect 3835 3488 4620 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4614 3476 4620 3488
rect 4672 3476 4678 3528
rect 5644 3525 5672 3692
rect 5902 3680 5908 3732
rect 5960 3680 5966 3732
rect 6270 3680 6276 3732
rect 6328 3680 6334 3732
rect 6730 3680 6736 3732
rect 6788 3680 6794 3732
rect 7650 3680 7656 3732
rect 7708 3680 7714 3732
rect 7006 3612 7012 3664
rect 7064 3652 7070 3664
rect 7837 3655 7895 3661
rect 7837 3652 7849 3655
rect 7064 3624 7849 3652
rect 7064 3612 7070 3624
rect 7837 3621 7849 3624
rect 7883 3621 7895 3655
rect 7837 3615 7895 3621
rect 6086 3544 6092 3596
rect 6144 3544 6150 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3584 6607 3587
rect 6595 3556 7420 3584
rect 6595 3553 6607 3556
rect 6549 3547 6607 3553
rect 5629 3519 5687 3525
rect 5629 3485 5641 3519
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 6362 3476 6368 3528
rect 6420 3476 6426 3528
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3516 7067 3519
rect 7282 3516 7288 3528
rect 7055 3488 7288 3516
rect 7055 3485 7067 3488
rect 7009 3479 7067 3485
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7392 3525 7420 3556
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 2222 3408 2228 3460
rect 2280 3408 2286 3460
rect 3142 3408 3148 3460
rect 3200 3448 3206 3460
rect 3237 3451 3295 3457
rect 3237 3448 3249 3451
rect 3200 3420 3249 3448
rect 3200 3408 3206 3420
rect 3237 3417 3249 3420
rect 3283 3417 3295 3451
rect 3237 3411 3295 3417
rect 6917 3451 6975 3457
rect 6917 3417 6929 3451
rect 6963 3448 6975 3451
rect 7098 3448 7104 3460
rect 6963 3420 7104 3448
rect 6963 3417 6975 3420
rect 6917 3411 6975 3417
rect 7098 3408 7104 3420
rect 7156 3408 7162 3460
rect 3418 3340 3424 3392
rect 3476 3389 3482 3392
rect 3476 3383 3495 3389
rect 3483 3349 3495 3383
rect 3476 3343 3495 3349
rect 3605 3383 3663 3389
rect 3605 3349 3617 3383
rect 3651 3380 3663 3383
rect 4706 3380 4712 3392
rect 3651 3352 4712 3380
rect 3651 3349 3663 3352
rect 3605 3343 3663 3349
rect 3476 3340 3482 3343
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 7282 3340 7288 3392
rect 7340 3380 7346 3392
rect 7392 3380 7420 3479
rect 8018 3476 8024 3528
rect 8076 3476 8082 3528
rect 7340 3352 7420 3380
rect 7340 3340 7346 3352
rect 7466 3340 7472 3392
rect 7524 3340 7530 3392
rect 1104 3290 8372 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 8372 3290
rect 1104 3216 8372 3238
rect 1026 3136 1032 3188
rect 1084 3176 1090 3188
rect 1489 3179 1547 3185
rect 1489 3176 1501 3179
rect 1084 3148 1501 3176
rect 1084 3136 1090 3148
rect 1489 3145 1501 3148
rect 1535 3145 1547 3179
rect 1489 3139 1547 3145
rect 2222 3136 2228 3188
rect 2280 3136 2286 3188
rect 3418 3136 3424 3188
rect 3476 3176 3482 3188
rect 3973 3179 4031 3185
rect 3973 3176 3985 3179
rect 3476 3148 3985 3176
rect 3476 3136 3482 3148
rect 3973 3145 3985 3148
rect 4019 3145 4031 3179
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 3973 3139 4031 3145
rect 4172 3148 6193 3176
rect 4062 3068 4068 3120
rect 4120 3108 4126 3120
rect 4172 3117 4200 3148
rect 6181 3145 6193 3148
rect 6227 3176 6239 3179
rect 6227 3148 6592 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 4157 3111 4215 3117
rect 4157 3108 4169 3111
rect 4120 3080 4169 3108
rect 4120 3068 4126 3080
rect 4157 3077 4169 3080
rect 4203 3077 4215 3111
rect 4157 3071 4215 3077
rect 4706 3068 4712 3120
rect 4764 3068 4770 3120
rect 6457 3111 6515 3117
rect 6457 3108 6469 3111
rect 5934 3080 6469 3108
rect 6457 3077 6469 3080
rect 6503 3077 6515 3111
rect 6457 3071 6515 3077
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 1673 3043 1731 3049
rect 1673 3040 1685 3043
rect 1452 3012 1685 3040
rect 1452 3000 1458 3012
rect 1673 3009 1685 3012
rect 1719 3009 1731 3043
rect 1673 3003 1731 3009
rect 2133 3043 2191 3049
rect 2133 3009 2145 3043
rect 2179 3040 2191 3043
rect 2406 3040 2412 3052
rect 2179 3012 2412 3040
rect 2179 3009 2191 3012
rect 2133 3003 2191 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 3786 3000 3792 3052
rect 3844 3040 3850 3052
rect 4341 3043 4399 3049
rect 4341 3040 4353 3043
rect 3844 3012 4353 3040
rect 3844 3000 3850 3012
rect 4341 3009 4353 3012
rect 4387 3009 4399 3043
rect 4341 3003 4399 3009
rect 4430 3000 4436 3052
rect 4488 3000 4494 3052
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 6564 2972 6592 3148
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 7377 3179 7435 3185
rect 7377 3176 7389 3179
rect 7156 3148 7389 3176
rect 7156 3136 7162 3148
rect 7377 3145 7389 3148
rect 7423 3145 7435 3179
rect 7377 3139 7435 3145
rect 7282 3068 7288 3120
rect 7340 3068 7346 3120
rect 6914 3000 6920 3052
rect 6972 3000 6978 3052
rect 7006 3000 7012 3052
rect 7064 3040 7070 3052
rect 7591 3043 7649 3049
rect 7591 3040 7603 3043
rect 7064 3012 7109 3040
rect 7208 3012 7603 3040
rect 7064 3000 7070 3012
rect 7208 2972 7236 3012
rect 7591 3009 7603 3012
rect 7637 3009 7649 3043
rect 7591 3003 7649 3009
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 7834 3040 7840 3052
rect 7791 3012 7840 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 8018 3000 8024 3052
rect 8076 3000 8082 3052
rect 6564 2944 7236 2972
rect 7024 2916 7052 2944
rect 7006 2864 7012 2916
rect 7064 2864 7070 2916
rect 7834 2796 7840 2848
rect 7892 2796 7898 2848
rect 1104 2746 8372 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 8372 2746
rect 1104 2672 8372 2694
rect 7466 2524 7472 2576
rect 7524 2524 7530 2576
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 7064 2400 7113 2428
rect 7064 2388 7070 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7255 2431 7313 2437
rect 7255 2397 7267 2431
rect 7301 2428 7313 2431
rect 7834 2428 7840 2440
rect 7301 2400 7840 2428
rect 7301 2397 7313 2400
rect 7255 2391 7313 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 1104 2202 8372 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 8372 2202
rect 1104 2128 8372 2150
<< via1 >>
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 4068 9120 4120 9172
rect 3792 9052 3844 9104
rect 3148 8848 3200 8900
rect 4804 8916 4856 8968
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 4068 8780 4120 8832
rect 4712 8780 4764 8832
rect 4804 8823 4856 8832
rect 4804 8789 4813 8823
rect 4813 8789 4847 8823
rect 4847 8789 4856 8823
rect 4804 8780 4856 8789
rect 6644 8780 6696 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 4620 8508 4672 8560
rect 5724 8508 5776 8560
rect 6644 8483 6696 8492
rect 6644 8449 6653 8483
rect 6653 8449 6687 8483
rect 6687 8449 6696 8483
rect 6644 8440 6696 8449
rect 3148 8372 3200 8424
rect 4804 8372 4856 8424
rect 6828 8440 6880 8492
rect 7472 8440 7524 8492
rect 6920 8304 6972 8356
rect 3148 8236 3200 8288
rect 3884 8236 3936 8288
rect 6092 8236 6144 8288
rect 6184 8279 6236 8288
rect 6184 8245 6193 8279
rect 6193 8245 6227 8279
rect 6227 8245 6236 8279
rect 6184 8236 6236 8245
rect 7380 8279 7432 8288
rect 7380 8245 7389 8279
rect 7389 8245 7423 8279
rect 7423 8245 7432 8279
rect 7380 8236 7432 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3056 8032 3108 8084
rect 3792 8032 3844 8084
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6000 8075 6052 8084
rect 6000 8041 6009 8075
rect 6009 8041 6043 8075
rect 6043 8041 6052 8075
rect 6000 8032 6052 8041
rect 6828 8032 6880 8084
rect 3884 8007 3936 8016
rect 3884 7973 3893 8007
rect 3893 7973 3927 8007
rect 3927 7973 3936 8007
rect 3884 7964 3936 7973
rect 4252 7964 4304 8016
rect 4896 7964 4948 8016
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 2228 7760 2280 7812
rect 2780 7692 2832 7744
rect 4712 7896 4764 7948
rect 4528 7828 4580 7880
rect 5080 7828 5132 7880
rect 6000 7896 6052 7948
rect 6092 7896 6144 7948
rect 5724 7828 5776 7880
rect 3424 7735 3476 7744
rect 3424 7701 3451 7735
rect 3451 7701 3476 7735
rect 3424 7692 3476 7701
rect 6184 7828 6236 7880
rect 7380 7896 7432 7948
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 7104 7760 7156 7812
rect 4160 7692 4212 7744
rect 4436 7692 4488 7744
rect 4528 7735 4580 7744
rect 4528 7701 4537 7735
rect 4537 7701 4571 7735
rect 4571 7701 4580 7735
rect 4528 7692 4580 7701
rect 4804 7692 4856 7744
rect 6736 7692 6788 7744
rect 6920 7735 6972 7744
rect 6920 7701 6929 7735
rect 6929 7701 6963 7735
rect 6963 7701 6972 7735
rect 6920 7692 6972 7701
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 2780 7420 2832 7472
rect 2412 7352 2464 7404
rect 2688 7395 2740 7404
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 3424 7420 3476 7472
rect 5264 7488 5316 7540
rect 7012 7488 7064 7540
rect 7472 7488 7524 7540
rect 4896 7420 4948 7472
rect 3792 7395 3844 7404
rect 3792 7361 3801 7395
rect 3801 7361 3835 7395
rect 3835 7361 3844 7395
rect 3792 7352 3844 7361
rect 4252 7395 4304 7404
rect 4252 7361 4265 7395
rect 4265 7361 4304 7395
rect 4252 7352 4304 7361
rect 4528 7352 4580 7404
rect 5264 7352 5316 7404
rect 6276 7352 6328 7404
rect 4344 7284 4396 7336
rect 4712 7284 4764 7336
rect 4160 7148 4212 7200
rect 4896 7216 4948 7268
rect 8024 7395 8076 7404
rect 8024 7361 8033 7395
rect 8033 7361 8067 7395
rect 8067 7361 8076 7395
rect 8024 7352 8076 7361
rect 4804 7148 4856 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 4804 6944 4856 6996
rect 3148 6851 3200 6860
rect 3148 6817 3157 6851
rect 3157 6817 3191 6851
rect 3191 6817 3200 6851
rect 3148 6808 3200 6817
rect 4896 6808 4948 6860
rect 6092 6808 6144 6860
rect 3332 6783 3384 6792
rect 3332 6749 3341 6783
rect 3341 6749 3375 6783
rect 3375 6749 3384 6783
rect 3332 6740 3384 6749
rect 2136 6672 2188 6724
rect 2872 6715 2924 6724
rect 2872 6681 2881 6715
rect 2881 6681 2915 6715
rect 2915 6681 2924 6715
rect 2872 6672 2924 6681
rect 2688 6604 2740 6656
rect 6644 6783 6696 6792
rect 6644 6749 6653 6783
rect 6653 6749 6687 6783
rect 6687 6749 6696 6783
rect 6644 6740 6696 6749
rect 6736 6783 6788 6792
rect 6736 6749 6745 6783
rect 6745 6749 6779 6783
rect 6779 6749 6788 6783
rect 6736 6740 6788 6749
rect 4712 6672 4764 6724
rect 5540 6672 5592 6724
rect 4160 6604 4212 6656
rect 4252 6647 4304 6656
rect 4252 6613 4261 6647
rect 4261 6613 4295 6647
rect 4295 6613 4304 6647
rect 4252 6604 4304 6613
rect 4896 6604 4948 6656
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2872 6400 2924 6452
rect 5540 6400 5592 6452
rect 2688 6332 2740 6384
rect 3056 6375 3108 6384
rect 3056 6341 3065 6375
rect 3065 6341 3099 6375
rect 3099 6341 3108 6375
rect 3056 6332 3108 6341
rect 4160 6332 4212 6384
rect 5172 6332 5224 6384
rect 5356 6332 5408 6384
rect 848 6264 900 6316
rect 2412 6264 2464 6316
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 7012 6264 7064 6316
rect 7104 6307 7156 6316
rect 7104 6273 7113 6307
rect 7113 6273 7147 6307
rect 7147 6273 7156 6307
rect 7104 6264 7156 6273
rect 7380 6307 7432 6316
rect 7380 6273 7389 6307
rect 7389 6273 7423 6307
rect 7423 6273 7432 6307
rect 7380 6264 7432 6273
rect 1768 6060 1820 6112
rect 2228 6060 2280 6112
rect 3332 6128 3384 6180
rect 3976 6060 4028 6112
rect 4252 6060 4304 6112
rect 4620 6060 4672 6112
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 6276 6128 6328 6180
rect 6920 6060 6972 6112
rect 7288 6060 7340 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 5356 5856 5408 5908
rect 6644 5899 6696 5908
rect 6644 5865 6653 5899
rect 6653 5865 6687 5899
rect 6687 5865 6696 5899
rect 6644 5856 6696 5865
rect 7288 5899 7340 5908
rect 7288 5865 7297 5899
rect 7297 5865 7331 5899
rect 7331 5865 7340 5899
rect 7288 5856 7340 5865
rect 7472 5899 7524 5908
rect 7472 5865 7481 5899
rect 7481 5865 7515 5899
rect 7515 5865 7524 5899
rect 7472 5856 7524 5865
rect 4804 5788 4856 5840
rect 6736 5788 6788 5840
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 4160 5720 4212 5772
rect 4896 5720 4948 5772
rect 2412 5652 2464 5704
rect 4068 5652 4120 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7012 5652 7064 5704
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 3332 5584 3384 5636
rect 4252 5584 4304 5636
rect 5264 5584 5316 5636
rect 7656 5584 7708 5636
rect 2780 5516 2832 5568
rect 3792 5516 3844 5568
rect 4712 5516 4764 5568
rect 6920 5516 6972 5568
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 3976 5312 4028 5364
rect 2044 5244 2096 5296
rect 2780 5244 2832 5296
rect 5264 5312 5316 5364
rect 5632 5244 5684 5296
rect 4160 5176 4212 5228
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7288 5312 7340 5364
rect 6920 5244 6972 5296
rect 3332 5040 3384 5092
rect 4252 5040 4304 5092
rect 3884 4972 3936 5024
rect 5356 5108 5408 5160
rect 7380 5176 7432 5228
rect 8024 5219 8076 5228
rect 8024 5185 8033 5219
rect 8033 5185 8067 5219
rect 8067 5185 8076 5219
rect 8024 5176 8076 5185
rect 7104 5108 7156 5160
rect 7564 5108 7616 5160
rect 4712 4972 4764 5024
rect 6920 4972 6972 5024
rect 7472 4972 7524 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 5632 4768 5684 4820
rect 7748 4811 7800 4820
rect 7748 4777 7757 4811
rect 7757 4777 7791 4811
rect 7791 4777 7800 4811
rect 7748 4768 7800 4777
rect 3792 4700 3844 4752
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 4068 4632 4120 4684
rect 7288 4632 7340 4684
rect 7564 4675 7616 4684
rect 7564 4641 7573 4675
rect 7573 4641 7607 4675
rect 7607 4641 7616 4675
rect 7564 4632 7616 4641
rect 4804 4564 4856 4616
rect 5540 4564 5592 4616
rect 6184 4564 6236 4616
rect 6920 4607 6972 4616
rect 6920 4573 6929 4607
rect 6929 4573 6963 4607
rect 6963 4573 6972 4607
rect 6920 4564 6972 4573
rect 7472 4607 7524 4616
rect 7472 4573 7481 4607
rect 7481 4573 7515 4607
rect 7515 4573 7524 4607
rect 7472 4564 7524 4573
rect 2228 4539 2280 4548
rect 2228 4505 2237 4539
rect 2237 4505 2271 4539
rect 2271 4505 2280 4539
rect 2228 4496 2280 4505
rect 3056 4496 3108 4548
rect 5356 4496 5408 4548
rect 6368 4471 6420 4480
rect 6368 4437 6377 4471
rect 6377 4437 6411 4471
rect 6411 4437 6420 4471
rect 6368 4428 6420 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 3792 4131 3844 4140
rect 3792 4097 3801 4131
rect 3801 4097 3835 4131
rect 3835 4097 3844 4131
rect 3792 4088 3844 4097
rect 4068 4088 4120 4140
rect 4712 4156 4764 4208
rect 6276 4156 6328 4208
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7012 4088 7064 4097
rect 1400 4020 1452 4072
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 5908 4020 5960 4072
rect 6920 4020 6972 4072
rect 2872 3927 2924 3936
rect 2872 3893 2881 3927
rect 2881 3893 2915 3927
rect 2915 3893 2924 3927
rect 2872 3884 2924 3893
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 5724 3884 5776 3936
rect 7288 3884 7340 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 1400 3723 1452 3732
rect 1400 3689 1409 3723
rect 1409 3689 1443 3723
rect 1443 3689 1452 3723
rect 1400 3680 1452 3689
rect 3884 3680 3936 3732
rect 2872 3587 2924 3596
rect 2872 3553 2881 3587
rect 2881 3553 2915 3587
rect 2915 3553 2924 3587
rect 2872 3544 2924 3553
rect 4436 3544 4488 3596
rect 4712 3544 4764 3596
rect 4620 3476 4672 3528
rect 5908 3723 5960 3732
rect 5908 3689 5917 3723
rect 5917 3689 5951 3723
rect 5951 3689 5960 3723
rect 5908 3680 5960 3689
rect 6276 3723 6328 3732
rect 6276 3689 6285 3723
rect 6285 3689 6319 3723
rect 6319 3689 6328 3723
rect 6276 3680 6328 3689
rect 6736 3723 6788 3732
rect 6736 3689 6745 3723
rect 6745 3689 6779 3723
rect 6779 3689 6788 3723
rect 6736 3680 6788 3689
rect 7656 3723 7708 3732
rect 7656 3689 7665 3723
rect 7665 3689 7699 3723
rect 7699 3689 7708 3723
rect 7656 3680 7708 3689
rect 7012 3612 7064 3664
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 6368 3519 6420 3528
rect 6368 3485 6377 3519
rect 6377 3485 6411 3519
rect 6411 3485 6420 3519
rect 6368 3476 6420 3485
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 2228 3408 2280 3460
rect 3148 3408 3200 3460
rect 7104 3451 7156 3460
rect 7104 3417 7113 3451
rect 7113 3417 7147 3451
rect 7147 3417 7156 3451
rect 7104 3408 7156 3417
rect 3424 3383 3476 3392
rect 3424 3349 3449 3383
rect 3449 3349 3476 3383
rect 3424 3340 3476 3349
rect 4712 3340 4764 3392
rect 7288 3340 7340 3392
rect 8024 3519 8076 3528
rect 8024 3485 8033 3519
rect 8033 3485 8067 3519
rect 8067 3485 8076 3519
rect 8024 3476 8076 3485
rect 7472 3383 7524 3392
rect 7472 3349 7481 3383
rect 7481 3349 7515 3383
rect 7515 3349 7524 3383
rect 7472 3340 7524 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1032 3136 1084 3188
rect 2228 3179 2280 3188
rect 2228 3145 2237 3179
rect 2237 3145 2271 3179
rect 2271 3145 2280 3179
rect 2228 3136 2280 3145
rect 3424 3136 3476 3188
rect 4068 3068 4120 3120
rect 4712 3111 4764 3120
rect 4712 3077 4721 3111
rect 4721 3077 4755 3111
rect 4755 3077 4764 3111
rect 4712 3068 4764 3077
rect 1400 3000 1452 3052
rect 2412 3000 2464 3052
rect 3792 3000 3844 3052
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7104 3136 7156 3188
rect 7288 3111 7340 3120
rect 7288 3077 7297 3111
rect 7297 3077 7331 3111
rect 7331 3077 7340 3111
rect 7288 3068 7340 3077
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 7012 3043 7064 3052
rect 7012 3009 7022 3043
rect 7022 3009 7056 3043
rect 7056 3009 7064 3043
rect 7012 3000 7064 3009
rect 7840 3000 7892 3052
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 7012 2864 7064 2916
rect 7840 2839 7892 2848
rect 7840 2805 7849 2839
rect 7849 2805 7883 2839
rect 7883 2805 7892 2839
rect 7840 2796 7892 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 7472 2567 7524 2576
rect 7472 2533 7481 2567
rect 7481 2533 7515 2567
rect 7515 2533 7524 2567
rect 7472 2524 7524 2533
rect 7012 2388 7064 2440
rect 7840 2388 7892 2440
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 3882 10962 3938 11629
rect 4526 10962 4582 11629
rect 6458 10962 6514 11629
rect 3882 10934 4108 10962
rect 3882 10829 3938 10934
rect 4080 9178 4108 10934
rect 4526 10934 4844 10962
rect 4526 10829 4582 10934
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 3160 8430 3188 8842
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3160 8294 3188 8366
rect 3148 8288 3200 8294
rect 3148 8230 3200 8236
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 2240 7546 2268 7754
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2792 7478 2820 7686
rect 3068 7546 3096 8026
rect 3160 7886 3188 8230
rect 3804 8090 3832 9046
rect 4816 8974 4844 10934
rect 6458 10934 6592 10962
rect 6458 10829 6514 10934
rect 6564 8974 6592 10934
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 846 6352 902 6361
rect 846 6287 848 6296
rect 900 6287 902 6296
rect 848 6258 900 6264
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1780 5710 1808 6054
rect 2148 5914 2176 6666
rect 2424 6322 2452 7346
rect 2700 6662 2728 7346
rect 3054 6896 3110 6905
rect 3160 6866 3188 7822
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3436 7478 3464 7686
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3804 7410 3832 8026
rect 3896 8022 3924 8230
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 4080 7886 4108 8774
rect 4620 8560 4672 8566
rect 4620 8502 4672 8508
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4252 8016 4304 8022
rect 4252 7958 4304 7964
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 4160 7744 4212 7750
rect 4160 7686 4212 7692
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 4172 7206 4200 7686
rect 4264 7410 4292 7958
rect 4528 7880 4580 7886
rect 4356 7828 4528 7834
rect 4356 7822 4580 7828
rect 4356 7806 4568 7822
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4356 7342 4384 7806
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4528 7744 4580 7750
rect 4528 7686 4580 7692
rect 4448 7546 4476 7686
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4540 7410 4568 7686
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4344 7336 4396 7342
rect 4344 7278 4396 7284
rect 4160 7200 4212 7206
rect 4160 7142 4212 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3054 6831 3110 6840
rect 3148 6860 3200 6866
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6390 2728 6598
rect 2884 6458 2912 6666
rect 2872 6452 2924 6458
rect 2872 6394 2924 6400
rect 3068 6390 3096 6831
rect 3148 6802 3200 6808
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 2044 5296 2096 5302
rect 2044 5238 2096 5244
rect 2056 4826 2084 5238
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2240 4554 2268 6054
rect 2424 5710 2452 6258
rect 3344 6186 3372 6734
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4172 6390 4200 6598
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2228 4548 2280 4554
rect 2228 4490 2280 4496
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1412 3738 1440 4014
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1030 3496 1086 3505
rect 1030 3431 1086 3440
rect 1044 3194 1072 3431
rect 1032 3188 1084 3194
rect 1032 3130 1084 3136
rect 1412 3058 1440 3674
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 2240 3194 2268 3402
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2424 3058 2452 5646
rect 3344 5642 3372 6122
rect 3976 6112 4028 6118
rect 4172 6100 4200 6326
rect 4264 6118 4292 6598
rect 4632 6118 4660 8502
rect 4724 7954 4752 8774
rect 4816 8514 4844 8774
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5724 8560 5776 8566
rect 4816 8486 4936 8514
rect 5724 8502 5776 8508
rect 4804 8424 4856 8430
rect 4804 8366 4856 8372
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4816 7834 4844 8366
rect 4908 8022 4936 8486
rect 5736 8090 5764 8502
rect 6656 8498 6684 8774
rect 6644 8492 6696 8498
rect 6644 8434 6696 8440
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 6012 7954 6040 8026
rect 6104 7954 6132 8230
rect 6000 7948 6052 7954
rect 6000 7890 6052 7896
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6196 7886 6224 8230
rect 6840 8090 6868 8434
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 4724 7806 4844 7834
rect 5080 7880 5132 7886
rect 5724 7880 5776 7886
rect 5132 7828 5304 7834
rect 5080 7822 5304 7828
rect 5724 7822 5776 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6932 7834 6960 8298
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7392 7954 7420 8230
rect 7380 7948 7432 7954
rect 7380 7890 7432 7896
rect 7484 7886 7512 8434
rect 7472 7880 7524 7886
rect 5092 7806 5304 7822
rect 4724 7342 4752 7806
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4816 7206 4844 7686
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 5276 7546 5304 7806
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 4896 7472 4948 7478
rect 4896 7414 4948 7420
rect 4908 7274 4936 7414
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4804 6996 4856 7002
rect 4804 6938 4856 6944
rect 4712 6724 4764 6730
rect 4712 6666 4764 6672
rect 3976 6054 4028 6060
rect 4080 6072 4200 6100
rect 4252 6112 4304 6118
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 2792 5302 2820 5510
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 3332 5092 3384 5098
rect 3332 5034 3384 5040
rect 3344 4622 3372 5034
rect 3804 4758 3832 5510
rect 3988 5370 4016 6054
rect 4080 5710 4108 6072
rect 4252 6054 4304 6060
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 4172 5234 4200 5714
rect 4252 5636 4304 5642
rect 4252 5578 4304 5584
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4172 5114 4200 5170
rect 4080 5086 4200 5114
rect 4264 5098 4292 5578
rect 4252 5092 4304 5098
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4826 3924 4966
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3792 4752 3844 4758
rect 3792 4694 3844 4700
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3068 4078 3096 4490
rect 3804 4146 3832 4694
rect 4080 4690 4108 5086
rect 4252 5034 4304 5040
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2884 3602 2912 3878
rect 2872 3596 2924 3602
rect 2872 3538 2924 3544
rect 3068 3448 3096 4014
rect 3148 3460 3200 3466
rect 3068 3420 3148 3448
rect 3148 3402 3200 3408
rect 3424 3392 3476 3398
rect 3424 3334 3476 3340
rect 3436 3194 3464 3334
rect 3424 3188 3476 3194
rect 3424 3130 3476 3136
rect 3804 3058 3832 4082
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3738 3924 3878
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 4080 3126 4108 4082
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4068 3120 4120 3126
rect 4068 3062 4120 3068
rect 4448 3058 4476 3538
rect 4632 3534 4660 6054
rect 4724 5574 4752 6666
rect 4816 5846 4844 6938
rect 4908 6866 4936 7210
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4908 6662 4936 6802
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5172 6384 5224 6390
rect 5276 6338 5304 7346
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5552 6458 5580 6666
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5224 6332 5304 6338
rect 5172 6326 5304 6332
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5184 6310 5304 6326
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4804 5840 4856 5846
rect 4804 5782 4856 5788
rect 4908 5778 4936 6054
rect 5368 5914 5396 6326
rect 5540 6316 5592 6322
rect 5736 6304 5764 7822
rect 6932 7818 7144 7834
rect 7472 7822 7524 7828
rect 6932 7812 7156 7818
rect 6932 7806 7104 7812
rect 6932 7750 6960 7806
rect 7104 7754 7156 7760
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6920 7744 6972 7750
rect 6920 7686 6972 7692
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6092 6860 6144 6866
rect 6092 6802 6144 6808
rect 5592 6276 5764 6304
rect 5540 6258 5592 6264
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 4896 5772 4948 5778
rect 4896 5714 4948 5720
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 4712 5568 4764 5574
rect 4764 5528 4844 5556
rect 4712 5510 4764 5516
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4214 4752 4966
rect 4816 4622 4844 5528
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5276 5370 5304 5578
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5368 5166 5396 5850
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 5368 4554 5396 5102
rect 5552 4622 5580 6258
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5644 4826 5672 5238
rect 5632 4820 5684 4826
rect 5632 4762 5684 4768
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4724 3602 4752 4150
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 5736 3534 5764 3878
rect 5920 3738 5948 4014
rect 5908 3732 5960 3738
rect 5908 3674 5960 3680
rect 6104 3602 6132 6802
rect 6288 6662 6316 7346
rect 6748 6798 6776 7686
rect 7024 7546 7052 7686
rect 7484 7546 7512 7822
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8036 6905 8064 7346
rect 8022 6896 8078 6905
rect 8022 6831 8078 6840
rect 6644 6792 6696 6798
rect 6644 6734 6696 6740
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6186 6316 6598
rect 6276 6180 6328 6186
rect 6276 6122 6328 6128
rect 6656 5914 6684 6734
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6736 5840 6788 5846
rect 6736 5782 6788 5788
rect 6184 4616 6236 4622
rect 6184 4558 6236 4564
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 4620 3528 4672 3534
rect 4620 3470 4672 3476
rect 5724 3528 5776 3534
rect 6196 3516 6224 4558
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6288 3738 6316 4150
rect 6380 4146 6408 4422
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6748 3738 6776 5782
rect 6932 5710 6960 6054
rect 7024 5710 7052 6258
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 6932 5302 6960 5510
rect 7024 5370 7052 5510
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 5296 6972 5302
rect 6920 5238 6972 5244
rect 6932 5030 6960 5238
rect 7116 5166 7144 6258
rect 7392 6225 7420 6258
rect 7378 6216 7434 6225
rect 7378 6151 7434 6160
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7300 5914 7328 6054
rect 7484 5914 7512 6734
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7300 5370 7328 5850
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7104 5160 7156 5166
rect 7104 5102 7156 5108
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 7300 4690 7328 5306
rect 7392 5234 7420 5646
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7484 4622 7512 4966
rect 7576 4690 7604 5102
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 7472 4616 7524 4622
rect 7472 4558 7524 4564
rect 6932 4078 6960 4558
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6276 3732 6328 3738
rect 6276 3674 6328 3680
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6368 3528 6420 3534
rect 6196 3488 6368 3516
rect 5724 3470 5776 3476
rect 6368 3470 6420 3476
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3126 4752 3334
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 6380 3058 6408 3470
rect 6932 3058 6960 4014
rect 7024 3670 7052 4082
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 7024 3058 7052 3606
rect 7300 3534 7328 3878
rect 7668 3738 7696 5578
rect 7760 4826 7788 5646
rect 8022 5536 8078 5545
rect 8022 5471 8078 5480
rect 8036 5234 8064 5471
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7288 3528 7340 3534
rect 8024 3528 8076 3534
rect 7288 3470 7340 3476
rect 8022 3496 8024 3505
rect 8076 3496 8078 3505
rect 7104 3460 7156 3466
rect 8022 3431 8078 3440
rect 7104 3402 7156 3408
rect 7116 3194 7144 3402
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7472 3392 7524 3398
rect 7472 3334 7524 3340
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7300 3126 7328 3334
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7012 2916 7064 2922
rect 7012 2858 7064 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 7024 2446 7052 2858
rect 7484 2582 7512 3334
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7852 2854 7880 2994
rect 7840 2848 7892 2854
rect 8036 2825 8064 2994
rect 7840 2790 7892 2796
rect 8022 2816 8078 2825
rect 7472 2576 7524 2582
rect 7472 2518 7524 2524
rect 7852 2446 7880 2790
rect 8022 2751 8078 2760
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
<< via2 >>
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 846 6316 902 6352
rect 846 6296 848 6316
rect 848 6296 900 6316
rect 900 6296 902 6316
rect 3054 6840 3110 6896
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 1030 3440 1086 3496
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 8022 6840 8078 6896
rect 7378 6160 7434 6216
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 8022 5480 8078 5536
rect 8022 3476 8024 3496
rect 8024 3476 8076 3496
rect 8076 3476 8078 3496
rect 8022 3440 8078 3476
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 8022 2760 8078 2816
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 0 6898 800 6928
rect 3049 6898 3115 6901
rect 0 6896 3115 6898
rect 0 6840 3054 6896
rect 3110 6840 3115 6896
rect 0 6838 3115 6840
rect 0 6808 800 6838
rect 3049 6835 3115 6838
rect 8017 6898 8083 6901
rect 8685 6898 9485 6928
rect 8017 6896 9485 6898
rect 8017 6840 8022 6896
rect 8078 6840 9485 6896
rect 8017 6838 9485 6840
rect 8017 6835 8083 6838
rect 8685 6808 9485 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 841 6354 907 6357
rect 798 6352 907 6354
rect 798 6296 846 6352
rect 902 6296 907 6352
rect 798 6291 907 6296
rect 798 6248 858 6291
rect 0 6158 858 6248
rect 7373 6218 7439 6221
rect 8685 6218 9485 6248
rect 7373 6216 9485 6218
rect 7373 6160 7378 6216
rect 7434 6160 9485 6216
rect 7373 6158 9485 6160
rect 0 6128 800 6158
rect 7373 6155 7439 6158
rect 8685 6128 9485 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 8017 5538 8083 5541
rect 8685 5538 9485 5568
rect 8017 5536 9485 5538
rect 8017 5480 8022 5536
rect 8078 5480 9485 5536
rect 8017 5478 9485 5480
rect 8017 5475 8083 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 8685 5448 9485 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 0 3498 800 3528
rect 1025 3498 1091 3501
rect 0 3496 1091 3498
rect 0 3440 1030 3496
rect 1086 3440 1091 3496
rect 0 3438 1091 3440
rect 0 3408 800 3438
rect 1025 3435 1091 3438
rect 8017 3498 8083 3501
rect 8685 3498 9485 3528
rect 8017 3496 9485 3498
rect 8017 3440 8022 3496
rect 8078 3440 9485 3496
rect 8017 3438 9485 3440
rect 8017 3435 8083 3438
rect 8685 3408 9485 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 8017 2818 8083 2821
rect 8685 2818 9485 2848
rect 8017 2816 9485 2818
rect 8017 2760 8022 2816
rect 8078 2760 9485 2816
rect 8017 2758 9485 2760
rect 8017 2755 8083 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 8685 2728 9485 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 9280 4528 9296
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 8736 5188 9296
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _056_
timestamp -25199
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _057_
timestamp -25199
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp -25199
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _059_
timestamp -25199
transform 1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp -25199
transform -1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _061_
timestamp -25199
transform -1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _062_
timestamp -25199
transform -1 0 4784 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _063_
timestamp -25199
transform 1 0 4048 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _064_
timestamp -25199
transform 1 0 3864 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _065_
timestamp -25199
transform 1 0 6624 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _066_
timestamp -25199
transform -1 0 7268 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _067_
timestamp -25199
transform -1 0 7820 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _068_
timestamp -25199
transform -1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _069_
timestamp -25199
transform -1 0 7544 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _070_
timestamp -25199
transform 1 0 6440 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _071_
timestamp -25199
transform -1 0 7820 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _072_
timestamp -25199
transform 1 0 6992 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _073_
timestamp -25199
transform 1 0 6900 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _074_
timestamp -25199
transform 1 0 7084 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _075_
timestamp -25199
transform 1 0 7084 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _076_
timestamp -25199
transform 1 0 6992 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _077_
timestamp -25199
transform -1 0 7820 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _078_
timestamp -25199
transform 1 0 6900 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _079_
timestamp -25199
transform 1 0 6624 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _080_
timestamp -25199
transform 1 0 6532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _081_
timestamp -25199
transform 1 0 7452 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _082_
timestamp -25199
transform -1 0 7544 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _083_
timestamp -25199
transform -1 0 3404 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _084_
timestamp -25199
transform 1 0 2300 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _085_
timestamp -25199
transform 1 0 2668 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _086_
timestamp -25199
transform -1 0 4048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _087_
timestamp -25199
transform -1 0 3680 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _088_
timestamp -25199
transform -1 0 4968 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _089_
timestamp -25199
transform 1 0 4968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _090_
timestamp -25199
transform -1 0 5152 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _091_
timestamp -25199
transform 1 0 3220 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _092_
timestamp -25199
transform 1 0 3956 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _093_
timestamp -25199
transform 1 0 3864 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _094_
timestamp -25199
transform -1 0 5336 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _095_
timestamp -25199
transform -1 0 4324 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _096_
timestamp -25199
transform 1 0 3680 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _097_
timestamp -25199
transform -1 0 4876 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _098_
timestamp -25199
transform -1 0 3588 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _099_
timestamp -25199
transform -1 0 2668 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp -25199
transform 1 0 3772 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _101_
timestamp -25199
transform -1 0 4416 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _102_
timestamp -25199
transform 1 0 3220 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _103_
timestamp -25199
transform -1 0 6164 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _104_
timestamp -25199
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _105_
timestamp -25199
transform -1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp -25199
transform 1 0 5520 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _107_
timestamp -25199
transform -1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp -25199
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp -25199
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _110_
timestamp -25199
transform -1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp -25199
transform 1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _112_
timestamp -25199
transform -1 0 3220 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _113_
timestamp -25199
transform -1 0 3220 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _114_
timestamp -25199
transform 1 0 4416 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _115_
timestamp -25199
transform 1 0 4508 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _116_
timestamp -25199
transform 1 0 4324 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _117_
timestamp -25199
transform 1 0 1472 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _118_
timestamp -25199
transform 1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _119_
timestamp -25199
transform 1 0 4416 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp -25199
transform -1 0 3220 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp -25199
transform 1 0 3036 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp -25199
transform 1 0 3772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp -25199
transform -1 0 4416 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp -25199
transform -1 0 3496 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636943256
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636943256
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp -25199
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636943256
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636943256
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp -25199
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp -25199
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70
timestamp -25199
transform 1 0 7544 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp -25199
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_14
timestamp 1636943256
transform 1 0 2392 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_26
timestamp -25199
transform 1 0 3496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_30
timestamp -25199
transform 1 0 3864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_60
timestamp -25199
transform 1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_58
timestamp -25199
transform 1 0 6440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp -25199
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp -25199
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_9
timestamp -25199
transform 1 0 1932 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp -25199
transform 1 0 3404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_32
timestamp -25199
transform 1 0 4048 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp -25199
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_69
timestamp -25199
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_75
timestamp -25199
transform 1 0 8004 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_3
timestamp -25199
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_9
timestamp -25199
transform 1 0 1932 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_17
timestamp -25199
transform 1 0 2668 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_21
timestamp -25199
transform 1 0 3036 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp -25199
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp -25199
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_35
timestamp 1636943256
transform 1 0 4324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_50
timestamp -25199
transform 1 0 5704 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_56
timestamp -25199
transform 1 0 6256 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_73
timestamp -25199
transform 1 0 7820 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp -25199
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp -25199
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp -25199
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_60
timestamp -25199
transform 1 0 6624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_72
timestamp -25199
transform 1 0 7728 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_9
timestamp -25199
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_16
timestamp 1636943256
transform 1 0 2576 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_29
timestamp -25199
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636943256
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_53
timestamp -25199
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp -25199
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp -25199
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_19
timestamp -25199
transform 1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_46
timestamp -25199
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp -25199
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp -25199
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_57
timestamp -25199
transform 1 0 6348 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_7_66
timestamp -25199
transform 1 0 7176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp -25199
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp -25199
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_70
timestamp -25199
transform 1 0 7544 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_3
timestamp -25199
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_14
timestamp -25199
transform 1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_22
timestamp -25199
transform 1 0 3128 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_28
timestamp -25199
transform 1 0 3680 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_44
timestamp 1636943256
transform 1 0 5152 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp -25199
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_61
timestamp -25199
transform 1 0 6716 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp -25199
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_36
timestamp -25199
transform 1 0 4416 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_45
timestamp -25199
transform 1 0 5244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_55
timestamp -25199
transform 1 0 6164 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_70
timestamp -25199
transform 1 0 7544 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636943256
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_15
timestamp -25199
transform 1 0 2484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp -25199
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_11_69
timestamp -25199
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_75
timestamp -25199
transform 1 0 8004 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636943256
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp -25199
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_19
timestamp -25199
transform 1 0 2852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp -25199
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_46
timestamp -25199
transform 1 0 5336 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp -25199
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp -25199
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_62
timestamp 1636943256
transform 1 0 6808 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_74
timestamp -25199
transform 1 0 7912 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp -25199
transform 1 0 2024 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp -25199
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp -25199
transform -1 0 7084 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp -25199
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp -25199
transform 1 0 5060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp -25199
transform -1 0 6808 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp -25199
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp -25199
transform -1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp -25199
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp -25199
transform 1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp -25199
transform 1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input9
timestamp -25199
transform -1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output10
timestamp -25199
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp -25199
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp -25199
transform -1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp -25199
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp -25199
transform -1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp -25199
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp -25199
transform -1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp -25199
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp -25199
transform -1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp -25199
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp -25199
transform -1 0 8372 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp -25199
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp -25199
transform -1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp -25199
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp -25199
transform -1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp -25199
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp -25199
transform -1 0 8372 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp -25199
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp -25199
transform -1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp -25199
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp -25199
transform -1 0 8372 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp -25199
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp -25199
transform -1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp -25199
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp -25199
transform -1 0 8372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp -25199
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp -25199
transform -1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26
timestamp -25199
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp -25199
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp -25199
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp -25199
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_30
timestamp -25199
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_31
timestamp -25199
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_32
timestamp -25199
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_33
timestamp -25199
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_34
timestamp -25199
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_35
timestamp -25199
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_36
timestamp -25199
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_37
timestamp -25199
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_38
timestamp -25199
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_39
timestamp -25199
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_40
timestamp -25199
transform 1 0 6256 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 out
port 3 nsew signal output
flabel metal2 s 4526 10829 4582 11629 0 FreeSans 224 90 0 0 psc[0]
port 4 nsew signal input
flabel metal2 s 3882 10829 3938 11629 0 FreeSans 224 90 0 0 psc[1]
port 5 nsew signal input
flabel metal2 s 6458 10829 6514 11629 0 FreeSans 224 90 0 0 psc[2]
port 6 nsew signal input
flabel metal3 s 8685 6808 9485 6928 0 FreeSans 480 0 0 0 psc[3]
port 7 nsew signal input
flabel metal3 s 8685 6128 9485 6248 0 FreeSans 480 0 0 0 psc[4]
port 8 nsew signal input
flabel metal3 s 8685 5448 9485 5568 0 FreeSans 480 0 0 0 psc[5]
port 9 nsew signal input
flabel metal3 s 8685 2728 9485 2848 0 FreeSans 480 0 0 0 psc[6]
port 10 nsew signal input
flabel metal3 s 8685 3408 9485 3528 0 FreeSans 480 0 0 0 psc[7]
port 11 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 rst
port 12 nsew signal input
rlabel metal1 4738 8704 4738 8704 0 VGND
rlabel metal1 4738 9248 4738 9248 0 VPWR
rlabel metal1 2852 6426 2852 6426 0 _000_
rlabel metal1 3082 7786 3082 7786 0 _001_
rlabel metal1 4554 7276 4554 7276 0 _002_
rlabel metal1 4738 6834 4738 6834 0 _003_
rlabel metal1 4646 5304 4646 5304 0 _004_
rlabel metal2 2070 5032 2070 5032 0 _005_
rlabel metal2 4738 3230 4738 3230 0 _006_
rlabel metal2 5934 3876 5934 3876 0 _007_
rlabel metal2 2162 6290 2162 6290 0 _008_
rlabel metal2 2254 7650 2254 7650 0 _009_
rlabel metal2 5750 8296 5750 8296 0 _010_
rlabel metal1 5612 6426 5612 6426 0 _011_
rlabel metal1 5612 4794 5612 4794 0 _012_
rlabel metal2 2806 5406 2806 5406 0 _013_
rlabel metal1 6217 3094 6217 3094 0 _014_
rlabel metal2 6302 3944 6302 3944 0 _015_
rlabel metal2 2254 3298 2254 3298 0 _016_
rlabel metal2 2898 3740 2898 3740 0 _017_
rlabel metal2 5750 3706 5750 3706 0 _018_
rlabel metal2 6946 5406 6946 5406 0 _019_
rlabel metal2 7314 5984 7314 5984 0 _020_
rlabel metal1 6440 8058 6440 8058 0 _021_
rlabel metal2 4094 8330 4094 8330 0 _022_
rlabel metal1 4232 7786 4232 7786 0 _023_
rlabel metal1 4416 7832 4416 7832 0 _024_
rlabel metal1 6532 7854 6532 7854 0 _025_
rlabel metal2 6946 8024 6946 8024 0 _026_
rlabel metal2 7038 7616 7038 7616 0 _027_
rlabel metal2 7498 8160 7498 8160 0 _028_
rlabel metal1 7268 7922 7268 7922 0 _029_
rlabel metal1 6785 7922 6785 7922 0 _030_
rlabel metal1 6624 7718 6624 7718 0 _031_
rlabel metal2 7130 3298 7130 3298 0 _032_
rlabel metal2 7314 3706 7314 3706 0 _033_
rlabel metal1 7406 3536 7406 3536 0 _034_
rlabel metal2 7498 2958 7498 2958 0 _035_
rlabel metal1 7866 5644 7866 5644 0 _036_
rlabel metal2 7038 5440 7038 5440 0 _037_
rlabel metal2 7774 5236 7774 5236 0 _038_
rlabel metal2 6946 5882 6946 5882 0 _039_
rlabel metal2 6670 6324 6670 6324 0 _040_
rlabel metal2 6762 4760 6762 4760 0 _041_
rlabel metal2 7498 6324 7498 6324 0 _042_
rlabel metal1 4600 6630 4600 6630 0 _043_
rlabel metal2 3082 7786 3082 7786 0 _044_
rlabel metal1 4232 7446 4232 7446 0 _045_
rlabel metal1 5144 6358 5144 6358 0 _046_
rlabel metal1 4784 7174 4784 7174 0 _047_
rlabel metal1 4684 5542 4684 5542 0 _048_
rlabel metal1 4600 5814 4600 5814 0 _049_
rlabel metal1 3956 5202 3956 5202 0 _050_
rlabel metal2 3910 4896 3910 4896 0 _051_
rlabel metal2 3818 4828 3818 4828 0 _052_
rlabel metal1 2714 4794 2714 4794 0 _053_
rlabel metal1 4554 3706 4554 3706 0 _054_
rlabel metal1 3726 3162 3726 3162 0 _055_
rlabel metal3 1878 6868 1878 6868 0 clk
rlabel metal1 4600 6086 4600 6086 0 clknet_0_clk
rlabel metal1 2944 5134 2944 5134 0 clknet_1_0__leaf_clk
rlabel metal1 3864 6834 3864 6834 0 clknet_1_1__leaf_clk
rlabel via1 4263 7378 4263 7378 0 net1
rlabel metal2 1426 3876 1426 3876 0 net10
rlabel metal1 2944 4114 2944 4114 0 net11
rlabel metal2 1794 5882 1794 5882 0 net12
rlabel metal2 6394 4284 6394 4284 0 net13
rlabel metal1 4692 8874 4692 8874 0 net2
rlabel metal2 6670 8636 6670 8636 0 net3
rlabel metal1 7682 7242 7682 7242 0 net4
rlabel metal1 7636 6290 7636 6290 0 net5
rlabel metal1 7406 5134 7406 5134 0 net6
rlabel metal2 7866 2618 7866 2618 0 net7
rlabel via1 7038 3026 7038 3026 0 net8
rlabel metal2 6394 3264 6394 3264 0 net9
rlabel metal1 1288 3162 1288 3162 0 out
rlabel metal1 4922 8942 4922 8942 0 psc[0]
rlabel metal1 5198 8942 5198 8942 0 psc[1]
rlabel metal2 6578 9945 6578 9945 0 psc[2]
rlabel metal3 8380 6868 8380 6868 0 psc[3]
rlabel metal2 7406 6239 7406 6239 0 psc[4]
rlabel metal2 8050 5355 8050 5355 0 psc[5]
rlabel metal2 8050 2907 8050 2907 0 psc[6]
rlabel via2 8050 3485 8050 3485 0 psc[7]
rlabel metal1 2530 6358 2530 6358 0 psc_cnt\[0\]
rlabel metal1 2852 7446 2852 7446 0 psc_cnt\[1\]
rlabel metal1 5934 7820 5934 7820 0 psc_cnt\[2\]
rlabel metal1 3772 5610 3772 5610 0 psc_cnt\[3\]
rlabel metal1 5014 5882 5014 5882 0 psc_cnt\[4\]
rlabel metal1 5060 5610 5060 5610 0 psc_cnt\[5\]
rlabel metal1 4140 3094 4140 3094 0 psc_cnt\[6\]
rlabel metal2 6946 3536 6946 3536 0 psc_cnt\[7\]
rlabel metal3 751 6188 751 6188 0 rst
<< properties >>
string FIXED_BBOX 0 0 9485 11629
<< end >>
