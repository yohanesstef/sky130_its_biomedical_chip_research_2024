VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO clk_int_div
  CLASS BLOCK ;
  FOREIGN clk_int_div ;
  ORIGIN 0.000 0.000 ;
  SIZE 74.945 BY 85.665 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 73.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 73.680 ;
    END
  END VPWR
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END clk_i
  PIN clk_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 81.665 48.670 85.665 ;
    END
  END clk_o
  PIN cycl_count_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END cycl_count_o[0]
  PIN cycl_count_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END cycl_count_o[1]
  PIN cycl_count_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END cycl_count_o[2]
  PIN cycl_count_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 70.945 23.840 74.945 24.440 ;
    END
  END cycl_count_o[3]
  PIN cycl_count_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 70.945 37.440 74.945 38.040 ;
    END
  END cycl_count_o[4]
  PIN cycl_count_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 70.945 40.840 74.945 41.440 ;
    END
  END cycl_count_o[5]
  PIN cycl_count_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 70.945 44.240 74.945 44.840 ;
    END
  END cycl_count_o[6]
  PIN cycl_count_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 70.945 47.640 74.945 48.240 ;
    END
  END cycl_count_o[7]
  PIN div_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END div_i[0]
  PIN div_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END div_i[1]
  PIN div_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END div_i[2]
  PIN div_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END div_i[3]
  PIN div_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END div_i[4]
  PIN div_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END div_i[5]
  PIN div_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END div_i[6]
  PIN div_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END div_i[7]
  PIN div_ready_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.336500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 81.665 29.350 85.665 ;
    END
  END div_ready_o
  PIN div_valid_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 81.665 32.570 85.665 ;
    END
  END div_valid_i
  PIN en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 81.665 35.790 85.665 ;
    END
  END en_i
  PIN rst_ni
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 70.945 20.440 74.945 21.040 ;
    END
  END rst_ni
  PIN test_mode_en_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 81.665 42.230 85.665 ;
    END
  END test_mode_en_i
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 69.190 73.630 ;
      LAYER li1 ;
        RECT 5.520 10.795 69.000 73.525 ;
      LAYER met1 ;
        RECT 4.210 10.640 69.000 73.680 ;
      LAYER met2 ;
        RECT 4.230 81.385 28.790 81.665 ;
        RECT 29.630 81.385 32.010 81.665 ;
        RECT 32.850 81.385 35.230 81.665 ;
        RECT 36.070 81.385 41.670 81.665 ;
        RECT 42.510 81.385 48.110 81.665 ;
        RECT 48.950 81.385 67.530 81.665 ;
        RECT 4.230 4.280 67.530 81.385 ;
        RECT 4.230 4.000 35.230 4.280 ;
        RECT 36.070 4.000 38.450 4.280 ;
        RECT 39.290 4.000 41.670 4.280 ;
        RECT 42.510 4.000 67.530 4.280 ;
      LAYER met3 ;
        RECT 3.990 65.640 70.945 73.605 ;
        RECT 4.400 64.240 70.945 65.640 ;
        RECT 3.990 58.840 70.945 64.240 ;
        RECT 4.400 57.440 70.945 58.840 ;
        RECT 3.990 48.640 70.945 57.440 ;
        RECT 3.990 47.240 70.545 48.640 ;
        RECT 3.990 45.240 70.945 47.240 ;
        RECT 4.400 43.840 70.545 45.240 ;
        RECT 3.990 41.840 70.945 43.840 ;
        RECT 4.400 40.440 70.545 41.840 ;
        RECT 3.990 38.440 70.945 40.440 ;
        RECT 4.400 37.040 70.545 38.440 ;
        RECT 3.990 35.040 70.945 37.040 ;
        RECT 4.400 33.640 70.945 35.040 ;
        RECT 3.990 31.640 70.945 33.640 ;
        RECT 4.400 30.240 70.945 31.640 ;
        RECT 3.990 28.240 70.945 30.240 ;
        RECT 4.400 26.840 70.945 28.240 ;
        RECT 3.990 24.840 70.945 26.840 ;
        RECT 4.400 23.440 70.545 24.840 ;
        RECT 3.990 21.440 70.945 23.440 ;
        RECT 3.990 20.040 70.545 21.440 ;
        RECT 3.990 10.715 70.945 20.040 ;
      LAYER met4 ;
        RECT 46.295 17.855 46.625 55.585 ;
  END
END clk_int_div
END LIBRARY

