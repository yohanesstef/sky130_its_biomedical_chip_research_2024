magic
tech sky130A
magscale 1 2
timestamp 1730474680
<< nwell >>
rect -214 -314 214 348
<< pmos >>
rect -120 -214 120 286
<< pdiff >>
rect -178 274 -120 286
rect -178 -202 -166 274
rect -132 -202 -120 274
rect -178 -214 -120 -202
rect 120 274 178 286
rect 120 -202 132 274
rect 166 -202 178 274
rect 120 -214 178 -202
<< pdiffc >>
rect -166 -202 -132 274
rect 132 -202 166 274
<< poly >>
rect -120 286 120 312
rect -120 -261 120 -214
rect -120 -295 -104 -261
rect 104 -295 120 -261
rect -120 -311 120 -295
<< polycont >>
rect -104 -295 104 -261
<< locali >>
rect -166 274 -132 290
rect -166 -218 -132 -202
rect 132 274 166 290
rect 132 -218 166 -202
rect -120 -295 -104 -261
rect 104 -295 120 -261
<< viali >>
rect -166 -202 -132 274
rect 132 -202 166 274
rect -104 -295 104 -261
<< metal1 >>
rect -172 274 -126 286
rect -172 -202 -166 274
rect -132 -202 -126 274
rect -172 -214 -126 -202
rect 126 274 172 286
rect 126 -202 132 274
rect 166 -202 172 274
rect 126 -214 172 -202
rect -116 -261 116 -255
rect -116 -295 -104 -261
rect 104 -295 116 -261
rect -116 -301 116 -295
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2.5 l 1.2 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
