magic
tech sky130A
magscale 1 2
timestamp 1730474680
<< error_p >>
rect -29 567 29 573
rect -29 533 -17 567
rect -29 527 29 533
rect -29 373 29 379
rect -29 339 -17 373
rect -29 333 29 339
rect -29 265 29 271
rect -29 231 -17 265
rect -29 225 29 231
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -231 29 -225
rect -29 -265 -17 -231
rect -29 -271 29 -265
rect -29 -339 29 -333
rect -29 -373 -17 -339
rect -29 -379 29 -373
rect -29 -533 29 -527
rect -29 -567 -17 -533
rect -29 -573 29 -567
<< pwell >>
rect -211 -705 211 705
<< nmos >>
rect -15 411 15 495
rect -15 109 15 193
rect -15 -193 15 -109
rect -15 -495 15 -411
<< ndiff >>
rect -73 483 -15 495
rect -73 423 -61 483
rect -27 423 -15 483
rect -73 411 -15 423
rect 15 483 73 495
rect 15 423 27 483
rect 61 423 73 483
rect 15 411 73 423
rect -73 181 -15 193
rect -73 121 -61 181
rect -27 121 -15 181
rect -73 109 -15 121
rect 15 181 73 193
rect 15 121 27 181
rect 61 121 73 181
rect 15 109 73 121
rect -73 -121 -15 -109
rect -73 -181 -61 -121
rect -27 -181 -15 -121
rect -73 -193 -15 -181
rect 15 -121 73 -109
rect 15 -181 27 -121
rect 61 -181 73 -121
rect 15 -193 73 -181
rect -73 -423 -15 -411
rect -73 -483 -61 -423
rect -27 -483 -15 -423
rect -73 -495 -15 -483
rect 15 -423 73 -411
rect 15 -483 27 -423
rect 61 -483 73 -423
rect 15 -495 73 -483
<< ndiffc >>
rect -61 423 -27 483
rect 27 423 61 483
rect -61 121 -27 181
rect 27 121 61 181
rect -61 -181 -27 -121
rect 27 -181 61 -121
rect -61 -483 -27 -423
rect 27 -483 61 -423
<< psubdiff >>
rect -175 635 -79 669
rect 79 635 175 669
rect -175 573 -141 635
rect 141 573 175 635
rect -175 -635 -141 -573
rect 141 -635 175 -573
rect -175 -669 -79 -635
rect 79 -669 175 -635
<< psubdiffcont >>
rect -79 635 79 669
rect -175 -573 -141 573
rect 141 -573 175 573
rect -79 -669 79 -635
<< poly >>
rect -33 567 33 583
rect -33 533 -17 567
rect 17 533 33 567
rect -33 517 33 533
rect -15 495 15 517
rect -15 389 15 411
rect -33 373 33 389
rect -33 339 -17 373
rect 17 339 33 373
rect -33 323 33 339
rect -33 265 33 281
rect -33 231 -17 265
rect 17 231 33 265
rect -33 215 33 231
rect -15 193 15 215
rect -15 87 15 109
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -109 15 -87
rect -15 -215 15 -193
rect -33 -231 33 -215
rect -33 -265 -17 -231
rect 17 -265 33 -231
rect -33 -281 33 -265
rect -33 -339 33 -323
rect -33 -373 -17 -339
rect 17 -373 33 -339
rect -33 -389 33 -373
rect -15 -411 15 -389
rect -15 -517 15 -495
rect -33 -533 33 -517
rect -33 -567 -17 -533
rect 17 -567 33 -533
rect -33 -583 33 -567
<< polycont >>
rect -17 533 17 567
rect -17 339 17 373
rect -17 231 17 265
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -265 17 -231
rect -17 -373 17 -339
rect -17 -567 17 -533
<< locali >>
rect -175 635 -79 669
rect 79 635 175 669
rect -175 573 -141 635
rect 141 573 175 635
rect -33 533 -17 567
rect 17 533 33 567
rect -61 483 -27 499
rect -61 407 -27 423
rect 27 483 61 499
rect 27 407 61 423
rect -33 339 -17 373
rect 17 339 33 373
rect -33 231 -17 265
rect 17 231 33 265
rect -61 181 -27 197
rect -61 105 -27 121
rect 27 181 61 197
rect 27 105 61 121
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -121 -27 -105
rect -61 -197 -27 -181
rect 27 -121 61 -105
rect 27 -197 61 -181
rect -33 -265 -17 -231
rect 17 -265 33 -231
rect -33 -373 -17 -339
rect 17 -373 33 -339
rect -61 -423 -27 -407
rect -61 -499 -27 -483
rect 27 -423 61 -407
rect 27 -499 61 -483
rect -33 -567 -17 -533
rect 17 -567 33 -533
rect -175 -635 -141 -573
rect 141 -635 175 -573
rect -175 -669 -79 -635
rect 79 -669 175 -635
<< viali >>
rect -17 533 17 567
rect -61 423 -27 483
rect 27 423 61 483
rect -17 339 17 373
rect -17 231 17 265
rect -61 121 -27 181
rect 27 121 61 181
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -181 -27 -121
rect 27 -181 61 -121
rect -17 -265 17 -231
rect -17 -373 17 -339
rect -61 -483 -27 -423
rect 27 -483 61 -423
rect -17 -567 17 -533
<< metal1 >>
rect -29 567 29 573
rect -29 533 -17 567
rect 17 533 29 567
rect -29 527 29 533
rect -67 483 -21 495
rect -67 423 -61 483
rect -27 423 -21 483
rect -67 411 -21 423
rect 21 483 67 495
rect 21 423 27 483
rect 61 423 67 483
rect 21 411 67 423
rect -29 373 29 379
rect -29 339 -17 373
rect 17 339 29 373
rect -29 333 29 339
rect -29 265 29 271
rect -29 231 -17 265
rect 17 231 29 265
rect -29 225 29 231
rect -67 181 -21 193
rect -67 121 -61 181
rect -27 121 -21 181
rect -67 109 -21 121
rect 21 181 67 193
rect 21 121 27 181
rect 61 121 67 181
rect 21 109 67 121
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -121 -21 -109
rect -67 -181 -61 -121
rect -27 -181 -21 -121
rect -67 -193 -21 -181
rect 21 -121 67 -109
rect 21 -181 27 -121
rect 61 -181 67 -121
rect 21 -193 67 -181
rect -29 -231 29 -225
rect -29 -265 -17 -231
rect 17 -265 29 -231
rect -29 -271 29 -265
rect -29 -339 29 -333
rect -29 -373 -17 -339
rect 17 -373 29 -339
rect -29 -379 29 -373
rect -67 -423 -21 -411
rect -67 -483 -61 -423
rect -27 -483 -21 -423
rect -67 -495 -21 -483
rect 21 -423 67 -411
rect 21 -483 27 -423
rect 61 -483 67 -423
rect 21 -495 67 -483
rect -29 -533 29 -527
rect -29 -567 -17 -533
rect 17 -567 29 -533
rect -29 -573 29 -567
<< properties >>
string FIXED_BBOX -158 -652 158 652
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.15 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
