magic
tech sky130A
magscale 1 2
timestamp 1729898924
<< checkpaint >>
rect -3932 -3932 16304 18448
<< viali >>
rect 8493 11849 8527 11883
rect 3985 11713 4019 11747
rect 4629 11713 4663 11747
rect 4905 11713 4939 11747
rect 5273 11713 5307 11747
rect 5917 11713 5951 11747
rect 7205 11713 7239 11747
rect 7849 11713 7883 11747
rect 8309 11713 8343 11747
rect 8401 11713 8435 11747
rect 8953 11713 8987 11747
rect 9229 11713 9263 11747
rect 8677 11645 8711 11679
rect 4169 11577 4203 11611
rect 4721 11577 4755 11611
rect 5457 11577 5491 11611
rect 7389 11577 7423 11611
rect 8033 11577 8067 11611
rect 4537 11509 4571 11543
rect 6101 11509 6135 11543
rect 8401 11509 8435 11543
rect 9137 11509 9171 11543
rect 9413 11509 9447 11543
rect 7941 11305 7975 11339
rect 8401 11305 8435 11339
rect 6193 11237 6227 11271
rect 8953 11169 8987 11203
rect 9321 11169 9355 11203
rect 10057 11169 10091 11203
rect 4353 11101 4387 11135
rect 5181 11101 5215 11135
rect 5365 11101 5399 11135
rect 5917 11101 5951 11135
rect 6101 11101 6135 11135
rect 6469 11101 6503 11135
rect 7205 11101 7239 11135
rect 7481 11101 7515 11135
rect 8032 11101 8066 11135
rect 8125 11101 8159 11135
rect 8492 11101 8526 11135
rect 8585 11101 8619 11135
rect 9413 11101 9447 11135
rect 9689 11101 9723 11135
rect 9843 11101 9877 11135
rect 4813 11033 4847 11067
rect 6193 11033 6227 11067
rect 7021 11033 7055 11067
rect 3801 10965 3835 10999
rect 6377 10965 6411 10999
rect 7389 10965 7423 10999
rect 9597 10965 9631 10999
rect 2881 10761 2915 10795
rect 3341 10693 3375 10727
rect 5917 10693 5951 10727
rect 2973 10625 3007 10659
rect 3433 10625 3467 10659
rect 3525 10625 3559 10659
rect 3985 10625 4019 10659
rect 4537 10625 4571 10659
rect 4721 10625 4755 10659
rect 5181 10625 5215 10659
rect 5273 10625 5307 10659
rect 5733 10625 5767 10659
rect 6101 10625 6135 10659
rect 7021 10625 7055 10659
rect 7389 10625 7423 10659
rect 8585 10625 8619 10659
rect 8677 10625 8711 10659
rect 8953 10625 8987 10659
rect 9045 10625 9079 10659
rect 9321 10625 9355 10659
rect 9414 10625 9448 10659
rect 9965 10625 9999 10659
rect 10057 10625 10091 10659
rect 2513 10557 2547 10591
rect 6653 10557 6687 10591
rect 6929 10557 6963 10591
rect 7573 10557 7607 10591
rect 7665 10557 7699 10591
rect 8033 10557 8067 10591
rect 9229 10557 9263 10591
rect 4353 10489 4387 10523
rect 8217 10489 8251 10523
rect 2697 10421 2731 10455
rect 3709 10421 3743 10455
rect 3893 10421 3927 10455
rect 8125 10421 8159 10455
rect 8769 10421 8803 10455
rect 9505 10421 9539 10455
rect 9781 10421 9815 10455
rect 3617 10217 3651 10251
rect 5089 10217 5123 10251
rect 6377 10217 6411 10251
rect 7941 10217 7975 10251
rect 8125 10217 8159 10251
rect 10885 10217 10919 10251
rect 4905 10149 4939 10183
rect 7205 10149 7239 10183
rect 7297 10149 7331 10183
rect 2145 10081 2179 10115
rect 4997 10081 5031 10115
rect 6193 10081 6227 10115
rect 9413 10081 9447 10115
rect 1869 10013 1903 10047
rect 4445 10013 4479 10047
rect 5457 10013 5491 10047
rect 5549 10013 5583 10047
rect 5733 10013 5767 10047
rect 5917 10013 5951 10047
rect 6009 10013 6043 10047
rect 6285 10013 6319 10047
rect 6561 10013 6595 10047
rect 7113 10013 7147 10047
rect 7389 10013 7423 10047
rect 7573 10013 7607 10047
rect 7757 10013 7791 10047
rect 8217 10013 8251 10047
rect 9137 10013 9171 10047
rect 6745 9945 6779 9979
rect 6929 9945 6963 9979
rect 3985 9877 4019 9911
rect 8217 9673 8251 9707
rect 9229 9673 9263 9707
rect 4077 9605 4111 9639
rect 8309 9605 8343 9639
rect 8493 9605 8527 9639
rect 10333 9605 10367 9639
rect 4721 9537 4755 9571
rect 4905 9537 4939 9571
rect 5181 9537 5215 9571
rect 5457 9537 5491 9571
rect 8125 9537 8159 9571
rect 8861 9537 8895 9571
rect 10241 9537 10275 9571
rect 2053 9469 2087 9503
rect 2329 9469 2363 9503
rect 5365 9469 5399 9503
rect 8953 9469 8987 9503
rect 3801 9401 3835 9435
rect 4445 9401 4479 9435
rect 5549 9401 5583 9435
rect 4537 9333 4571 9367
rect 7941 9333 7975 9367
rect 2789 9129 2823 9163
rect 2973 9129 3007 9163
rect 3893 9129 3927 9163
rect 4445 9129 4479 9163
rect 5365 9129 5399 9163
rect 5825 9129 5859 9163
rect 5181 9061 5215 9095
rect 6469 8993 6503 9027
rect 8309 8993 8343 9027
rect 8493 8993 8527 9027
rect 9045 8993 9079 9027
rect 3341 8925 3375 8959
rect 3525 8925 3559 8959
rect 4261 8925 4295 8959
rect 4537 8925 4571 8959
rect 6101 8925 6135 8959
rect 6377 8925 6411 8959
rect 6561 8925 6595 8959
rect 7297 8925 7331 8959
rect 8217 8925 8251 8959
rect 8401 8925 8435 8959
rect 2957 8857 2991 8891
rect 3157 8857 3191 8891
rect 4077 8857 4111 8891
rect 5349 8857 5383 8891
rect 5549 8857 5583 8891
rect 6009 8857 6043 8891
rect 7665 8857 7699 8891
rect 9321 8857 9355 8891
rect 3341 8789 3375 8823
rect 5641 8789 5675 8823
rect 5804 8789 5838 8823
rect 6193 8789 6227 8823
rect 8033 8789 8067 8823
rect 10793 8789 10827 8823
rect 4997 8585 5031 8619
rect 9045 8585 9079 8619
rect 9229 8585 9263 8619
rect 9689 8585 9723 8619
rect 10333 8585 10367 8619
rect 4629 8517 4663 8551
rect 1685 8449 1719 8483
rect 4905 8449 4939 8483
rect 5181 8449 5215 8483
rect 5365 8449 5399 8483
rect 6101 8449 6135 8483
rect 6377 8449 6411 8483
rect 6837 8449 6871 8483
rect 9321 8449 9355 8483
rect 9505 8449 9539 8483
rect 9597 8459 9631 8493
rect 9781 8449 9815 8483
rect 10241 8449 10275 8483
rect 2881 8381 2915 8415
rect 5549 8381 5583 8415
rect 7113 8381 7147 8415
rect 1501 8313 1535 8347
rect 4813 8313 4847 8347
rect 8585 8313 8619 8347
rect 8677 8313 8711 8347
rect 9321 8313 9355 8347
rect 6469 8245 6503 8279
rect 9045 8245 9079 8279
rect 3157 8041 3191 8075
rect 6745 8041 6779 8075
rect 7205 8041 7239 8075
rect 7665 8041 7699 8075
rect 7941 8041 7975 8075
rect 4629 7973 4663 8007
rect 6837 7973 6871 8007
rect 7389 7973 7423 8007
rect 3249 7905 3283 7939
rect 3893 7905 3927 7939
rect 4997 7905 5031 7939
rect 5273 7905 5307 7939
rect 1409 7837 1443 7871
rect 3433 7837 3467 7871
rect 4445 7837 4479 7871
rect 4629 7837 4663 7871
rect 4905 7837 4939 7871
rect 7757 7837 7791 7871
rect 7849 7837 7883 7871
rect 1685 7769 1719 7803
rect 7205 7769 7239 7803
rect 3617 7701 3651 7735
rect 4813 7701 4847 7735
rect 3341 7497 3375 7531
rect 5365 7497 5399 7531
rect 9321 7497 9355 7531
rect 8033 7429 8067 7463
rect 1777 7361 1811 7395
rect 2513 7361 2547 7395
rect 3157 7361 3191 7395
rect 3433 7361 3467 7395
rect 3617 7361 3651 7395
rect 5733 7361 5767 7395
rect 7849 7361 7883 7395
rect 1869 7293 1903 7327
rect 3893 7293 3927 7327
rect 1409 7225 1443 7259
rect 5825 7157 5859 7191
rect 6653 6953 6687 6987
rect 7389 6953 7423 6987
rect 1777 6817 1811 6851
rect 8953 6817 8987 6851
rect 3985 6749 4019 6783
rect 5365 6749 5399 6783
rect 7757 6749 7791 6783
rect 8033 6749 8067 6783
rect 2053 6681 2087 6715
rect 3893 6681 3927 6715
rect 9229 6681 9263 6715
rect 3525 6613 3559 6647
rect 7205 6613 7239 6647
rect 7389 6613 7423 6647
rect 7941 6613 7975 6647
rect 10701 6613 10735 6647
rect 2145 6409 2179 6443
rect 8493 6409 8527 6443
rect 8861 6409 8895 6443
rect 9505 6409 9539 6443
rect 10149 6409 10183 6443
rect 2605 6341 2639 6375
rect 5885 6341 5919 6375
rect 6101 6341 6135 6375
rect 7941 6341 7975 6375
rect 9321 6341 9355 6375
rect 9965 6341 9999 6375
rect 2697 6273 2731 6307
rect 5273 6273 5307 6307
rect 5457 6273 5491 6307
rect 8217 6273 8251 6307
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 8677 6273 8711 6307
rect 9597 6273 9631 6307
rect 9781 6273 9815 6307
rect 10241 6273 10275 6307
rect 2973 6205 3007 6239
rect 2329 6137 2363 6171
rect 5641 6137 5675 6171
rect 8953 6137 8987 6171
rect 4445 6069 4479 6103
rect 5733 6069 5767 6103
rect 5917 6069 5951 6103
rect 6469 6069 6503 6103
rect 9321 6069 9355 6103
rect 3065 5865 3099 5899
rect 3249 5865 3283 5899
rect 3893 5865 3927 5899
rect 4629 5865 4663 5899
rect 7205 5865 7239 5899
rect 7665 5865 7699 5899
rect 8125 5865 8159 5899
rect 8677 5865 8711 5899
rect 9137 5865 9171 5899
rect 10333 5865 10367 5899
rect 2973 5797 3007 5831
rect 4813 5729 4847 5763
rect 5089 5729 5123 5763
rect 7297 5729 7331 5763
rect 2329 5661 2363 5695
rect 2513 5661 2547 5695
rect 2789 5661 2823 5695
rect 3985 5661 4019 5695
rect 4537 5661 4571 5695
rect 4721 5661 4755 5695
rect 6745 5661 6779 5695
rect 7021 5661 7055 5695
rect 7481 5661 7515 5695
rect 7757 5661 7791 5695
rect 7941 5661 7975 5695
rect 8493 5661 8527 5695
rect 8677 5661 8711 5695
rect 9965 5661 9999 5695
rect 2605 5593 2639 5627
rect 3217 5593 3251 5627
rect 3433 5593 3467 5627
rect 8953 5593 8987 5627
rect 10609 5593 10643 5627
rect 2513 5525 2547 5559
rect 6561 5525 6595 5559
rect 6837 5525 6871 5559
rect 9153 5525 9187 5559
rect 9321 5525 9355 5559
rect 10057 5525 10091 5559
rect 2313 5321 2347 5355
rect 2605 5321 2639 5355
rect 4261 5321 4295 5355
rect 4537 5321 4571 5355
rect 7941 5321 7975 5355
rect 8401 5321 8435 5355
rect 2513 5253 2547 5287
rect 5549 5253 5583 5287
rect 8861 5253 8895 5287
rect 2605 5185 2639 5219
rect 2697 5185 2731 5219
rect 2881 5185 2915 5219
rect 4445 5185 4479 5219
rect 4629 5185 4663 5219
rect 5825 5185 5859 5219
rect 7757 5185 7791 5219
rect 7941 5185 7975 5219
rect 8217 5185 8251 5219
rect 8493 5185 8527 5219
rect 9137 5185 9171 5219
rect 8033 5117 8067 5151
rect 9413 5117 9447 5151
rect 4813 5049 4847 5083
rect 9045 5049 9079 5083
rect 2145 4981 2179 5015
rect 2329 4981 2363 5015
rect 8861 4981 8895 5015
rect 10885 4981 10919 5015
rect 3249 4777 3283 4811
rect 8585 4777 8619 4811
rect 1501 4641 1535 4675
rect 4353 4641 4387 4675
rect 8953 4641 8987 4675
rect 9229 4641 9263 4675
rect 3525 4573 3559 4607
rect 6377 4573 6411 4607
rect 8217 4573 8251 4607
rect 1777 4505 1811 4539
rect 3433 4505 3467 4539
rect 4629 4505 4663 4539
rect 6285 4505 6319 4539
rect 8401 4505 8435 4539
rect 6101 4437 6135 4471
rect 10701 4437 10735 4471
rect 2421 4233 2455 4267
rect 2789 4233 2823 4267
rect 4629 4233 4663 4267
rect 4905 4233 4939 4267
rect 8861 4233 8895 4267
rect 10701 4233 10735 4267
rect 6837 4165 6871 4199
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 4261 4097 4295 4131
rect 5181 4097 5215 4131
rect 5273 4097 5307 4131
rect 5365 4097 5399 4131
rect 6561 4097 6595 4131
rect 6653 4097 6687 4131
rect 7205 4097 7239 4131
rect 7389 4097 7423 4131
rect 7481 4097 7515 4131
rect 8309 4097 8343 4131
rect 8677 4097 8711 4131
rect 8861 4097 8895 4131
rect 9045 4097 9079 4131
rect 9137 4097 9171 4131
rect 10149 4097 10183 4131
rect 10241 4097 10275 4131
rect 10885 4097 10919 4131
rect 5089 4029 5123 4063
rect 7021 4029 7055 4063
rect 4813 3961 4847 3995
rect 4629 3893 4663 3927
rect 6837 3893 6871 3927
rect 8217 3893 8251 3927
rect 3893 3689 3927 3723
rect 5549 3689 5583 3723
rect 6837 3689 6871 3723
rect 7665 3689 7699 3723
rect 8125 3689 8159 3723
rect 8309 3621 8343 3655
rect 4353 3553 4387 3587
rect 6009 3553 6043 3587
rect 3801 3485 3835 3519
rect 4077 3485 4111 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 4813 3485 4847 3519
rect 5089 3485 5123 3519
rect 5365 3485 5399 3519
rect 5733 3485 5767 3519
rect 5917 3485 5951 3519
rect 6101 3485 6135 3519
rect 6285 3485 6319 3519
rect 7113 3485 7147 3519
rect 7849 3485 7883 3519
rect 7941 3485 7975 3519
rect 8217 3485 8251 3519
rect 8584 3485 8618 3519
rect 8677 3485 8711 3519
rect 4629 3417 4663 3451
rect 4721 3417 4755 3451
rect 6469 3417 6503 3451
rect 7389 3417 7423 3451
rect 4997 3349 5031 3383
rect 5181 3349 5215 3383
rect 7021 3349 7055 3383
rect 7205 3349 7239 3383
rect 4353 3145 4387 3179
rect 6469 3145 6503 3179
rect 7849 3145 7883 3179
rect 3617 3077 3651 3111
rect 4905 3077 4939 3111
rect 7481 3077 7515 3111
rect 8401 3077 8435 3111
rect 3525 3009 3559 3043
rect 3801 3009 3835 3043
rect 3893 3009 3927 3043
rect 4077 3009 4111 3043
rect 4169 3009 4203 3043
rect 4537 3009 4571 3043
rect 4813 3009 4847 3043
rect 5181 3009 5215 3043
rect 5273 3009 5307 3043
rect 6377 3009 6411 3043
rect 7020 3009 7054 3043
rect 7113 3009 7147 3043
rect 7205 3009 7239 3043
rect 7298 3009 7332 3043
rect 7573 3009 7607 3043
rect 7711 3009 7745 3043
rect 4629 2873 4663 2907
rect 7941 2873 7975 2907
rect 8125 2873 8159 2907
rect 6929 2805 6963 2839
rect 3525 2601 3559 2635
rect 4629 2601 4663 2635
rect 5273 2601 5307 2635
rect 6193 2601 6227 2635
rect 7297 2601 7331 2635
rect 8033 2601 8067 2635
rect 8677 2601 8711 2635
rect 4169 2533 4203 2567
rect 7389 2533 7423 2567
rect 6929 2465 6963 2499
rect 3341 2397 3375 2431
rect 3985 2397 4019 2431
rect 4813 2397 4847 2431
rect 5457 2397 5491 2431
rect 6009 2397 6043 2431
rect 6377 2397 6411 2431
rect 6531 2397 6565 2431
rect 6745 2397 6779 2431
rect 7113 2397 7147 2431
rect 7389 2397 7423 2431
rect 7573 2397 7607 2431
rect 7665 2397 7699 2431
rect 7757 2397 7791 2431
rect 8217 2397 8251 2431
rect 8493 2397 8527 2431
rect 7941 2261 7975 2295
<< metal1 >>
rect 1104 11994 11224 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 11224 11994
rect 1104 11920 11224 11942
rect 8481 11883 8539 11889
rect 8481 11849 8493 11883
rect 8527 11880 8539 11883
rect 9398 11880 9404 11892
rect 8527 11852 9404 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 4522 11772 4528 11824
rect 4580 11812 4586 11824
rect 4580 11784 4936 11812
rect 4580 11772 4586 11784
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4908 11753 4936 11784
rect 3973 11747 4031 11753
rect 3973 11744 3985 11747
rect 3936 11716 3985 11744
rect 3936 11704 3942 11716
rect 3973 11713 3985 11716
rect 4019 11713 4031 11747
rect 3973 11707 4031 11713
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11744 4675 11747
rect 4893 11747 4951 11753
rect 4663 11716 4752 11744
rect 4663 11713 4675 11716
rect 4617 11707 4675 11713
rect 4157 11611 4215 11617
rect 4157 11577 4169 11611
rect 4203 11608 4215 11611
rect 4614 11608 4620 11620
rect 4203 11580 4620 11608
rect 4203 11577 4215 11580
rect 4157 11571 4215 11577
rect 4614 11568 4620 11580
rect 4672 11568 4678 11620
rect 4724 11617 4752 11716
rect 4893 11713 4905 11747
rect 4939 11713 4951 11747
rect 4893 11707 4951 11713
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 5810 11704 5816 11756
rect 5868 11744 5874 11756
rect 5905 11747 5963 11753
rect 5905 11744 5917 11747
rect 5868 11716 5917 11744
rect 5868 11704 5874 11716
rect 5905 11713 5917 11716
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 7098 11704 7104 11756
rect 7156 11744 7162 11756
rect 7193 11747 7251 11753
rect 7193 11744 7205 11747
rect 7156 11716 7205 11744
rect 7156 11704 7162 11716
rect 7193 11713 7205 11716
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 7742 11704 7748 11756
rect 7800 11744 7806 11756
rect 7837 11747 7895 11753
rect 7837 11744 7849 11747
rect 7800 11716 7849 11744
rect 7800 11704 7806 11716
rect 7837 11713 7849 11716
rect 7883 11713 7895 11747
rect 7837 11707 7895 11713
rect 7926 11704 7932 11756
rect 7984 11744 7990 11756
rect 8297 11747 8355 11753
rect 8297 11744 8309 11747
rect 7984 11716 8309 11744
rect 7984 11704 7990 11716
rect 8297 11713 8309 11716
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8386 11704 8392 11756
rect 8444 11704 8450 11756
rect 8478 11704 8484 11756
rect 8536 11744 8542 11756
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8536 11716 8953 11744
rect 8536 11704 8542 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 9217 11747 9275 11753
rect 9217 11744 9229 11747
rect 9088 11716 9229 11744
rect 9088 11704 9094 11716
rect 9217 11713 9229 11716
rect 9263 11713 9275 11747
rect 9217 11707 9275 11713
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 9122 11676 9128 11688
rect 8711 11648 9128 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 9122 11636 9128 11648
rect 9180 11636 9186 11688
rect 4709 11611 4767 11617
rect 4709 11577 4721 11611
rect 4755 11577 4767 11611
rect 4709 11571 4767 11577
rect 5445 11611 5503 11617
rect 5445 11577 5457 11611
rect 5491 11608 5503 11611
rect 6454 11608 6460 11620
rect 5491 11580 6460 11608
rect 5491 11577 5503 11580
rect 5445 11571 5503 11577
rect 6454 11568 6460 11580
rect 6512 11568 6518 11620
rect 7377 11611 7435 11617
rect 7377 11577 7389 11611
rect 7423 11608 7435 11611
rect 7558 11608 7564 11620
rect 7423 11580 7564 11608
rect 7423 11577 7435 11580
rect 7377 11571 7435 11577
rect 7558 11568 7564 11580
rect 7616 11568 7622 11620
rect 8021 11611 8079 11617
rect 8021 11577 8033 11611
rect 8067 11608 8079 11611
rect 8294 11608 8300 11620
rect 8067 11580 8300 11608
rect 8067 11577 8079 11580
rect 8021 11571 8079 11577
rect 8294 11568 8300 11580
rect 8352 11608 8358 11620
rect 8938 11608 8944 11620
rect 8352 11580 8944 11608
rect 8352 11568 8358 11580
rect 8938 11568 8944 11580
rect 8996 11568 9002 11620
rect 4525 11543 4583 11549
rect 4525 11509 4537 11543
rect 4571 11540 4583 11543
rect 5166 11540 5172 11552
rect 4571 11512 5172 11540
rect 4571 11509 4583 11512
rect 4525 11503 4583 11509
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 6089 11543 6147 11549
rect 6089 11509 6101 11543
rect 6135 11540 6147 11543
rect 6270 11540 6276 11552
rect 6135 11512 6276 11540
rect 6135 11509 6147 11512
rect 6089 11503 6147 11509
rect 6270 11500 6276 11512
rect 6328 11500 6334 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 8389 11543 8447 11549
rect 8389 11540 8401 11543
rect 7524 11512 8401 11540
rect 7524 11500 7530 11512
rect 8389 11509 8401 11512
rect 8435 11509 8447 11543
rect 8389 11503 8447 11509
rect 8478 11500 8484 11552
rect 8536 11540 8542 11552
rect 9125 11543 9183 11549
rect 9125 11540 9137 11543
rect 8536 11512 9137 11540
rect 8536 11500 8542 11512
rect 9125 11509 9137 11512
rect 9171 11540 9183 11543
rect 9306 11540 9312 11552
rect 9171 11512 9312 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9401 11543 9459 11549
rect 9401 11509 9413 11543
rect 9447 11540 9459 11543
rect 9490 11540 9496 11552
rect 9447 11512 9496 11540
rect 9447 11509 9459 11512
rect 9401 11503 9459 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 1104 11450 11224 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 11224 11450
rect 1104 11376 11224 11398
rect 7926 11296 7932 11348
rect 7984 11296 7990 11348
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 5810 11228 5816 11280
rect 5868 11268 5874 11280
rect 6181 11271 6239 11277
rect 6181 11268 6193 11271
rect 5868 11240 6193 11268
rect 5868 11228 5874 11240
rect 6181 11237 6193 11240
rect 6227 11237 6239 11271
rect 6181 11231 6239 11237
rect 8294 11200 8300 11212
rect 7484 11172 8300 11200
rect 4338 11092 4344 11144
rect 4396 11092 4402 11144
rect 5166 11092 5172 11144
rect 5224 11092 5230 11144
rect 5350 11092 5356 11144
rect 5408 11092 5414 11144
rect 5905 11135 5963 11141
rect 5905 11101 5917 11135
rect 5951 11132 5963 11135
rect 5994 11132 6000 11144
rect 5951 11104 6000 11132
rect 5951 11101 5963 11104
rect 5905 11095 5963 11101
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6270 11132 6276 11144
rect 6135 11104 6276 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6270 11092 6276 11104
rect 6328 11092 6334 11144
rect 6454 11092 6460 11144
rect 6512 11092 6518 11144
rect 7193 11135 7251 11141
rect 7193 11101 7205 11135
rect 7239 11132 7251 11135
rect 7374 11132 7380 11144
rect 7239 11104 7380 11132
rect 7239 11101 7251 11104
rect 7193 11095 7251 11101
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7484 11141 7512 11172
rect 8294 11160 8300 11172
rect 8352 11160 8358 11212
rect 8404 11200 8432 11296
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 8404 11172 8953 11200
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 9122 11160 9128 11212
rect 9180 11200 9186 11212
rect 9309 11203 9367 11209
rect 9309 11200 9321 11203
rect 9180 11172 9321 11200
rect 9180 11160 9186 11172
rect 9309 11169 9321 11172
rect 9355 11200 9367 11203
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9355 11172 10057 11200
rect 9355 11169 9367 11172
rect 9309 11163 9367 11169
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10045 11163 10103 11169
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 8020 11135 8078 11141
rect 8020 11101 8032 11135
rect 8066 11101 8078 11135
rect 8020 11095 8078 11101
rect 4798 11024 4804 11076
rect 4856 11024 4862 11076
rect 5626 11024 5632 11076
rect 5684 11064 5690 11076
rect 6181 11067 6239 11073
rect 6181 11064 6193 11067
rect 5684 11036 6193 11064
rect 5684 11024 5690 11036
rect 6181 11033 6193 11036
rect 6227 11033 6239 11067
rect 6181 11027 6239 11033
rect 7009 11067 7067 11073
rect 7009 11033 7021 11067
rect 7055 11064 7067 11067
rect 7834 11064 7840 11076
rect 7055 11036 7840 11064
rect 7055 11033 7067 11036
rect 7009 11027 7067 11033
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 8036 11064 8064 11095
rect 8110 11092 8116 11144
rect 8168 11092 8174 11144
rect 8478 11132 8484 11144
rect 8439 11104 8484 11132
rect 8478 11092 8484 11104
rect 8536 11092 8542 11144
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 9214 11132 9220 11144
rect 8628 11104 9220 11132
rect 8628 11092 8634 11104
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9858 11141 9864 11144
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 9831 11135 9864 11141
rect 9831 11101 9843 11135
rect 9916 11132 9922 11144
rect 10870 11132 10876 11144
rect 9916 11104 10876 11132
rect 9831 11095 9864 11101
rect 9490 11064 9496 11076
rect 8036 11036 9496 11064
rect 9490 11024 9496 11036
rect 9548 11064 9554 11076
rect 9692 11064 9720 11095
rect 9858 11092 9864 11095
rect 9916 11092 9922 11104
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 9548 11036 9720 11064
rect 9548 11024 9554 11036
rect 3786 10956 3792 11008
rect 3844 10956 3850 11008
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6365 10999 6423 11005
rect 6365 10996 6377 10999
rect 5960 10968 6377 10996
rect 5960 10956 5966 10968
rect 6365 10965 6377 10968
rect 6411 10965 6423 10999
rect 6365 10959 6423 10965
rect 7377 10999 7435 11005
rect 7377 10965 7389 10999
rect 7423 10996 7435 10999
rect 7650 10996 7656 11008
rect 7423 10968 7656 10996
rect 7423 10965 7435 10968
rect 7377 10959 7435 10965
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 8294 10956 8300 11008
rect 8352 10996 8358 11008
rect 9585 10999 9643 11005
rect 9585 10996 9597 10999
rect 8352 10968 9597 10996
rect 8352 10956 8358 10968
rect 9585 10965 9597 10968
rect 9631 10965 9643 10999
rect 9585 10959 9643 10965
rect 1104 10906 11224 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 11224 10906
rect 1104 10832 11224 10854
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3786 10792 3792 10804
rect 2915 10764 3792 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7708 10764 9076 10792
rect 7708 10752 7714 10764
rect 3329 10727 3387 10733
rect 3329 10693 3341 10727
rect 3375 10724 3387 10727
rect 4338 10724 4344 10736
rect 3375 10696 4344 10724
rect 3375 10693 3387 10696
rect 3329 10687 3387 10693
rect 4338 10684 4344 10696
rect 4396 10724 4402 10736
rect 4396 10696 4752 10724
rect 4396 10684 4402 10696
rect 2958 10616 2964 10668
rect 3016 10616 3022 10668
rect 3421 10659 3479 10665
rect 3421 10625 3433 10659
rect 3467 10656 3479 10659
rect 3510 10656 3516 10668
rect 3467 10628 3516 10656
rect 3467 10625 3479 10628
rect 3421 10619 3479 10625
rect 3510 10616 3516 10628
rect 3568 10616 3574 10668
rect 3786 10616 3792 10668
rect 3844 10656 3850 10668
rect 3973 10659 4031 10665
rect 3973 10656 3985 10659
rect 3844 10628 3985 10656
rect 3844 10616 3850 10628
rect 3973 10625 3985 10628
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 4614 10656 4620 10668
rect 4571 10628 4620 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 4724 10665 4752 10696
rect 5626 10684 5632 10736
rect 5684 10724 5690 10736
rect 5905 10727 5963 10733
rect 5905 10724 5917 10727
rect 5684 10696 5917 10724
rect 5684 10684 5690 10696
rect 5905 10693 5917 10696
rect 5951 10693 5963 10727
rect 5905 10687 5963 10693
rect 7558 10684 7564 10736
rect 7616 10724 7622 10736
rect 7616 10696 8708 10724
rect 7616 10684 7622 10696
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 5166 10616 5172 10668
rect 5224 10616 5230 10668
rect 5261 10659 5319 10665
rect 5261 10625 5273 10659
rect 5307 10656 5319 10659
rect 5350 10656 5356 10668
rect 5307 10628 5356 10656
rect 5307 10625 5319 10628
rect 5261 10619 5319 10625
rect 5350 10616 5356 10628
rect 5408 10616 5414 10668
rect 5718 10616 5724 10668
rect 5776 10616 5782 10668
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10656 6147 10659
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 6135 10628 7021 10656
rect 6135 10625 6147 10628
rect 6089 10619 6147 10625
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7377 10659 7435 10665
rect 7377 10656 7389 10659
rect 7340 10628 7389 10656
rect 7340 10616 7346 10628
rect 7377 10625 7389 10628
rect 7423 10625 7435 10659
rect 7377 10619 7435 10625
rect 7742 10616 7748 10668
rect 7800 10656 7806 10668
rect 8680 10665 8708 10696
rect 8573 10659 8631 10665
rect 8573 10656 8585 10659
rect 7800 10628 8585 10656
rect 7800 10616 7806 10628
rect 8573 10625 8585 10628
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 8665 10659 8723 10665
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 2501 10591 2559 10597
rect 2501 10557 2513 10591
rect 2547 10588 2559 10591
rect 2682 10588 2688 10600
rect 2547 10560 2688 10588
rect 2547 10557 2559 10560
rect 2501 10551 2559 10557
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 6641 10591 6699 10597
rect 6641 10557 6653 10591
rect 6687 10588 6699 10591
rect 6822 10588 6828 10600
rect 6687 10560 6828 10588
rect 6687 10557 6699 10560
rect 6641 10551 6699 10557
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 6914 10548 6920 10600
rect 6972 10548 6978 10600
rect 7561 10591 7619 10597
rect 7561 10557 7573 10591
rect 7607 10588 7619 10591
rect 7653 10591 7711 10597
rect 7653 10588 7665 10591
rect 7607 10560 7665 10588
rect 7607 10557 7619 10560
rect 7561 10551 7619 10557
rect 7653 10557 7665 10560
rect 7699 10557 7711 10591
rect 7653 10551 7711 10557
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 8021 10591 8079 10597
rect 8021 10588 8033 10591
rect 7892 10560 8033 10588
rect 7892 10548 7898 10560
rect 8021 10557 8033 10560
rect 8067 10557 8079 10591
rect 8588 10588 8616 10619
rect 8938 10616 8944 10668
rect 8996 10616 9002 10668
rect 9048 10665 9076 10764
rect 9214 10684 9220 10736
rect 9272 10724 9278 10736
rect 9272 10696 9444 10724
rect 9272 10684 9278 10696
rect 9033 10659 9091 10665
rect 9033 10625 9045 10659
rect 9079 10625 9091 10659
rect 9033 10619 9091 10625
rect 9306 10616 9312 10668
rect 9364 10616 9370 10668
rect 9416 10665 9444 10696
rect 9402 10659 9460 10665
rect 9402 10625 9414 10659
rect 9448 10625 9460 10659
rect 9402 10619 9460 10625
rect 9582 10616 9588 10668
rect 9640 10656 9646 10668
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9640 10628 9965 10656
rect 9640 10616 9646 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10042 10616 10048 10668
rect 10100 10616 10106 10668
rect 9217 10591 9275 10597
rect 9217 10588 9229 10591
rect 8588 10560 9229 10588
rect 8021 10551 8079 10557
rect 9217 10557 9229 10560
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 4341 10523 4399 10529
rect 4341 10489 4353 10523
rect 4387 10520 4399 10523
rect 5074 10520 5080 10532
rect 4387 10492 5080 10520
rect 4387 10489 4399 10492
rect 4341 10483 4399 10489
rect 5074 10480 5080 10492
rect 5132 10480 5138 10532
rect 7926 10480 7932 10532
rect 7984 10520 7990 10532
rect 8205 10523 8263 10529
rect 8205 10520 8217 10523
rect 7984 10492 8217 10520
rect 7984 10480 7990 10492
rect 8205 10489 8217 10492
rect 8251 10489 8263 10523
rect 8205 10483 8263 10489
rect 2130 10412 2136 10464
rect 2188 10452 2194 10464
rect 2685 10455 2743 10461
rect 2685 10452 2697 10455
rect 2188 10424 2697 10452
rect 2188 10412 2194 10424
rect 2685 10421 2697 10424
rect 2731 10421 2743 10455
rect 2685 10415 2743 10421
rect 3694 10412 3700 10464
rect 3752 10412 3758 10464
rect 3878 10412 3884 10464
rect 3936 10412 3942 10464
rect 6546 10412 6552 10464
rect 6604 10452 6610 10464
rect 8113 10455 8171 10461
rect 8113 10452 8125 10455
rect 6604 10424 8125 10452
rect 6604 10412 6610 10424
rect 8113 10421 8125 10424
rect 8159 10421 8171 10455
rect 8113 10415 8171 10421
rect 8754 10412 8760 10464
rect 8812 10412 8818 10464
rect 9398 10412 9404 10464
rect 9456 10452 9462 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 9456 10424 9505 10452
rect 9456 10412 9462 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 9766 10412 9772 10464
rect 9824 10412 9830 10464
rect 1104 10362 11224 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 11224 10362
rect 1104 10288 11224 10310
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 3568 10220 3617 10248
rect 3568 10208 3574 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 3605 10211 3663 10217
rect 5074 10208 5080 10260
rect 5132 10208 5138 10260
rect 6365 10251 6423 10257
rect 6365 10217 6377 10251
rect 6411 10248 6423 10251
rect 6914 10248 6920 10260
rect 6411 10220 6920 10248
rect 6411 10217 6423 10220
rect 6365 10211 6423 10217
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 7374 10248 7380 10260
rect 7208 10220 7380 10248
rect 4893 10183 4951 10189
rect 4893 10149 4905 10183
rect 4939 10180 4951 10183
rect 6546 10180 6552 10192
rect 4939 10152 6552 10180
rect 4939 10149 4951 10152
rect 4893 10143 4951 10149
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 7208 10189 7236 10220
rect 7374 10208 7380 10220
rect 7432 10208 7438 10260
rect 7926 10208 7932 10260
rect 7984 10208 7990 10260
rect 8113 10251 8171 10257
rect 8113 10217 8125 10251
rect 8159 10248 8171 10251
rect 8754 10248 8760 10260
rect 8159 10220 8760 10248
rect 8159 10217 8171 10220
rect 8113 10211 8171 10217
rect 7193 10183 7251 10189
rect 7193 10149 7205 10183
rect 7239 10149 7251 10183
rect 7193 10143 7251 10149
rect 7285 10183 7343 10189
rect 7285 10149 7297 10183
rect 7331 10180 7343 10183
rect 7742 10180 7748 10192
rect 7331 10152 7748 10180
rect 7331 10149 7343 10152
rect 7285 10143 7343 10149
rect 7742 10140 7748 10152
rect 7800 10140 7806 10192
rect 2130 10072 2136 10124
rect 2188 10072 2194 10124
rect 4798 10072 4804 10124
rect 4856 10112 4862 10124
rect 4985 10115 5043 10121
rect 4985 10112 4997 10115
rect 4856 10084 4997 10112
rect 4856 10072 4862 10084
rect 4985 10081 4997 10084
rect 5031 10081 5043 10115
rect 5810 10112 5816 10124
rect 4985 10075 5043 10081
rect 5460 10084 5816 10112
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 1872 9976 1900 10007
rect 4154 10004 4160 10056
rect 4212 10044 4218 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 4212 10016 4445 10044
rect 4212 10004 4218 10016
rect 4433 10013 4445 10016
rect 4479 10044 4491 10047
rect 5350 10044 5356 10056
rect 4479 10016 5356 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 5460 10053 5488 10084
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 6178 10072 6184 10124
rect 6236 10072 6242 10124
rect 7944 10112 7972 10208
rect 7116 10084 7972 10112
rect 5445 10047 5503 10053
rect 5445 10013 5457 10047
rect 5491 10013 5503 10047
rect 5445 10007 5503 10013
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 5592 10016 5733 10044
rect 5592 10004 5598 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 5902 10004 5908 10056
rect 5960 10004 5966 10056
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 2038 9976 2044 9988
rect 1872 9948 2044 9976
rect 2038 9936 2044 9948
rect 2096 9936 2102 9988
rect 3878 9976 3884 9988
rect 3358 9948 3884 9976
rect 3878 9936 3884 9948
rect 3936 9936 3942 9988
rect 6012 9976 6040 10007
rect 6270 10004 6276 10056
rect 6328 10004 6334 10056
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 7116 10053 7144 10084
rect 7101 10047 7159 10053
rect 7101 10013 7113 10047
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 7377 10047 7435 10053
rect 7377 10013 7389 10047
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 6454 9976 6460 9988
rect 6012 9948 6460 9976
rect 6454 9936 6460 9948
rect 6512 9936 6518 9988
rect 6733 9979 6791 9985
rect 6733 9945 6745 9979
rect 6779 9976 6791 9979
rect 6917 9979 6975 9985
rect 6917 9976 6929 9979
rect 6779 9948 6929 9976
rect 6779 9945 6791 9948
rect 6733 9939 6791 9945
rect 6917 9945 6929 9948
rect 6963 9945 6975 9979
rect 7392 9976 7420 10007
rect 7558 10004 7564 10056
rect 7616 10004 7622 10056
rect 7745 10047 7803 10053
rect 7745 10013 7757 10047
rect 7791 10044 7803 10047
rect 8128 10044 8156 10211
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 10870 10208 10876 10260
rect 10928 10208 10934 10260
rect 9401 10115 9459 10121
rect 9401 10081 9413 10115
rect 9447 10112 9459 10115
rect 9766 10112 9772 10124
rect 9447 10084 9772 10112
rect 9447 10081 9459 10084
rect 9401 10075 9459 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 7791 10016 8156 10044
rect 7791 10013 7803 10016
rect 7745 10007 7803 10013
rect 8202 10004 8208 10056
rect 8260 10004 8266 10056
rect 9030 10004 9036 10056
rect 9088 10044 9094 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 9088 10016 9137 10044
rect 9088 10004 9094 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 8294 9976 8300 9988
rect 7392 9948 8300 9976
rect 6917 9939 6975 9945
rect 8294 9936 8300 9948
rect 8352 9936 8358 9988
rect 10410 9936 10416 9988
rect 10468 9936 10474 9988
rect 3970 9868 3976 9920
rect 4028 9868 4034 9920
rect 1104 9818 11224 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 11224 9818
rect 1104 9744 11224 9766
rect 8110 9664 8116 9716
rect 8168 9664 8174 9716
rect 8202 9664 8208 9716
rect 8260 9664 8266 9716
rect 9217 9707 9275 9713
rect 9217 9673 9229 9707
rect 9263 9704 9275 9707
rect 9582 9704 9588 9716
rect 9263 9676 9588 9704
rect 9263 9673 9275 9676
rect 9217 9667 9275 9673
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 3694 9596 3700 9648
rect 3752 9636 3758 9648
rect 4065 9639 4123 9645
rect 4065 9636 4077 9639
rect 3752 9608 4077 9636
rect 3752 9596 3758 9608
rect 4065 9605 4077 9608
rect 4111 9605 4123 9639
rect 5534 9636 5540 9648
rect 4065 9599 4123 9605
rect 4908 9608 5540 9636
rect 4709 9571 4767 9577
rect 2038 9460 2044 9512
rect 2096 9460 2102 9512
rect 2317 9503 2375 9509
rect 2317 9469 2329 9503
rect 2363 9500 2375 9503
rect 2774 9500 2780 9512
rect 2363 9472 2780 9500
rect 2363 9469 2375 9472
rect 2317 9463 2375 9469
rect 2774 9460 2780 9472
rect 2832 9460 2838 9512
rect 3436 9500 3464 9554
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 4798 9568 4804 9580
rect 4755 9540 4804 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 4908 9577 4936 9608
rect 5534 9596 5540 9608
rect 5592 9596 5598 9648
rect 8128 9636 8156 9664
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 8128 9608 8309 9636
rect 8297 9605 8309 9608
rect 8343 9605 8355 9639
rect 8297 9599 8355 9605
rect 8481 9639 8539 9645
rect 8481 9605 8493 9639
rect 8527 9636 8539 9639
rect 8570 9636 8576 9648
rect 8527 9608 8576 9636
rect 8527 9605 8539 9608
rect 8481 9599 8539 9605
rect 4893 9571 4951 9577
rect 4893 9537 4905 9571
rect 4939 9537 4951 9571
rect 4893 9531 4951 9537
rect 5169 9571 5227 9577
rect 5169 9537 5181 9571
rect 5215 9568 5227 9571
rect 5258 9568 5264 9580
rect 5215 9540 5264 9568
rect 5215 9537 5227 9540
rect 5169 9531 5227 9537
rect 5258 9528 5264 9540
rect 5316 9528 5322 9580
rect 5445 9571 5503 9577
rect 5445 9537 5457 9571
rect 5491 9568 5503 9571
rect 5810 9568 5816 9580
rect 5491 9540 5816 9568
rect 5491 9537 5503 9540
rect 5445 9531 5503 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 8110 9528 8116 9580
rect 8168 9528 8174 9580
rect 8312 9568 8340 9599
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 10321 9639 10379 9645
rect 10321 9605 10333 9639
rect 10367 9636 10379 9639
rect 10410 9636 10416 9648
rect 10367 9608 10416 9636
rect 10367 9605 10379 9608
rect 10321 9599 10379 9605
rect 10410 9596 10416 9608
rect 10468 9596 10474 9648
rect 8386 9568 8392 9580
rect 8312 9540 8392 9568
rect 8386 9528 8392 9540
rect 8444 9568 8450 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8444 9540 8861 9568
rect 8444 9528 8450 9540
rect 8849 9537 8861 9540
rect 8895 9568 8907 9571
rect 9858 9568 9864 9580
rect 8895 9540 9864 9568
rect 8895 9537 8907 9540
rect 8849 9531 8907 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 4062 9500 4068 9512
rect 3436 9472 4068 9500
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 5353 9503 5411 9509
rect 5353 9469 5365 9503
rect 5399 9500 5411 9503
rect 5718 9500 5724 9512
rect 5399 9472 5724 9500
rect 5399 9469 5411 9472
rect 5353 9463 5411 9469
rect 5718 9460 5724 9472
rect 5776 9460 5782 9512
rect 8941 9503 8999 9509
rect 8941 9469 8953 9503
rect 8987 9500 8999 9503
rect 9122 9500 9128 9512
rect 8987 9472 9128 9500
rect 8987 9469 8999 9472
rect 8941 9463 8999 9469
rect 9122 9460 9128 9472
rect 9180 9460 9186 9512
rect 3789 9435 3847 9441
rect 3789 9401 3801 9435
rect 3835 9432 3847 9435
rect 3878 9432 3884 9444
rect 3835 9404 3884 9432
rect 3835 9401 3847 9404
rect 3789 9395 3847 9401
rect 3878 9392 3884 9404
rect 3936 9432 3942 9444
rect 4154 9432 4160 9444
rect 3936 9404 4160 9432
rect 3936 9392 3942 9404
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 4433 9435 4491 9441
rect 4433 9401 4445 9435
rect 4479 9432 4491 9435
rect 4614 9432 4620 9444
rect 4479 9404 4620 9432
rect 4479 9401 4491 9404
rect 4433 9395 4491 9401
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 5537 9435 5595 9441
rect 5537 9401 5549 9435
rect 5583 9432 5595 9435
rect 5902 9432 5908 9444
rect 5583 9404 5908 9432
rect 5583 9401 5595 9404
rect 5537 9395 5595 9401
rect 5902 9392 5908 9404
rect 5960 9392 5966 9444
rect 4525 9367 4583 9373
rect 4525 9333 4537 9367
rect 4571 9364 4583 9367
rect 5626 9364 5632 9376
rect 4571 9336 5632 9364
rect 4571 9333 4583 9336
rect 4525 9327 4583 9333
rect 5626 9324 5632 9336
rect 5684 9324 5690 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 7929 9367 7987 9373
rect 7929 9364 7941 9367
rect 6604 9336 7941 9364
rect 6604 9324 6610 9336
rect 7929 9333 7941 9336
rect 7975 9333 7987 9367
rect 7929 9327 7987 9333
rect 1104 9274 11224 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 11224 9274
rect 1104 9200 11224 9222
rect 2774 9120 2780 9172
rect 2832 9120 2838 9172
rect 2961 9163 3019 9169
rect 2961 9129 2973 9163
rect 3007 9160 3019 9163
rect 3881 9163 3939 9169
rect 3881 9160 3893 9163
rect 3007 9132 3893 9160
rect 3007 9129 3019 9132
rect 2961 9123 3019 9129
rect 3881 9129 3893 9132
rect 3927 9129 3939 9163
rect 3881 9123 3939 9129
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4433 9163 4491 9169
rect 4433 9160 4445 9163
rect 4120 9132 4445 9160
rect 4120 9120 4126 9132
rect 4433 9129 4445 9132
rect 4479 9129 4491 9163
rect 4433 9123 4491 9129
rect 5353 9163 5411 9169
rect 5353 9129 5365 9163
rect 5399 9160 5411 9163
rect 5442 9160 5448 9172
rect 5399 9132 5448 9160
rect 5399 9129 5411 9132
rect 5353 9123 5411 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 5810 9120 5816 9172
rect 5868 9160 5874 9172
rect 6362 9160 6368 9172
rect 5868 9132 6368 9160
rect 5868 9120 5874 9132
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 3786 9052 3792 9104
rect 3844 9092 3850 9104
rect 5169 9095 5227 9101
rect 3844 9064 4476 9092
rect 3844 9052 3850 9064
rect 3970 9024 3976 9036
rect 3344 8996 3976 9024
rect 3344 8965 3372 8996
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8956 3571 8959
rect 4249 8959 4307 8965
rect 4249 8956 4261 8959
rect 3559 8928 4261 8956
rect 3559 8925 3571 8928
rect 3513 8919 3571 8925
rect 4249 8925 4261 8928
rect 4295 8956 4307 8959
rect 4338 8956 4344 8968
rect 4295 8928 4344 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4448 8956 4476 9064
rect 5169 9061 5181 9095
rect 5215 9092 5227 9095
rect 5258 9092 5264 9104
rect 5215 9064 5264 9092
rect 5215 9061 5227 9064
rect 5169 9055 5227 9061
rect 5258 9052 5264 9064
rect 5316 9052 5322 9104
rect 5534 9092 5540 9104
rect 5368 9064 5540 9092
rect 5368 9024 5396 9064
rect 5534 9052 5540 9064
rect 5592 9052 5598 9104
rect 8202 9052 8208 9104
rect 8260 9092 8266 9104
rect 8260 9064 9168 9092
rect 8260 9052 8266 9064
rect 8312 9033 8340 9064
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 4724 8996 5396 9024
rect 5552 8996 6469 9024
rect 4522 8956 4528 8968
rect 4448 8928 4528 8956
rect 4522 8916 4528 8928
rect 4580 8916 4586 8968
rect 2958 8897 2964 8900
rect 2945 8891 2964 8897
rect 2945 8857 2957 8891
rect 2945 8851 2964 8857
rect 2958 8848 2964 8851
rect 3016 8848 3022 8900
rect 3145 8891 3203 8897
rect 3145 8857 3157 8891
rect 3191 8888 3203 8891
rect 3191 8860 4016 8888
rect 3191 8857 3203 8860
rect 3145 8851 3203 8857
rect 2976 8820 3004 8848
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 2976 8792 3341 8820
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3988 8820 4016 8860
rect 4062 8848 4068 8900
rect 4120 8848 4126 8900
rect 4724 8888 4752 8996
rect 5552 8958 5580 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 8297 9027 8355 9033
rect 8297 8993 8309 9027
rect 8343 9024 8355 9027
rect 8481 9027 8539 9033
rect 8343 8996 8377 9024
rect 8343 8993 8355 8996
rect 8297 8987 8355 8993
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 8570 9024 8576 9036
rect 8527 8996 8576 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 9030 8984 9036 9036
rect 9088 8984 9094 9036
rect 9140 9024 9168 9064
rect 9398 9024 9404 9036
rect 9140 8996 9404 9024
rect 9398 8984 9404 8996
rect 9456 9024 9462 9036
rect 9950 9024 9956 9036
rect 9456 8996 9956 9024
rect 9456 8984 9462 8996
rect 9950 8984 9956 8996
rect 10008 8984 10014 9036
rect 5368 8930 5580 8958
rect 6089 8959 6147 8965
rect 6089 8956 6101 8959
rect 4356 8860 4752 8888
rect 4356 8820 4384 8860
rect 4798 8848 4804 8900
rect 4856 8888 4862 8900
rect 5368 8897 5396 8930
rect 6012 8928 6101 8956
rect 6012 8900 6040 8928
rect 6089 8925 6101 8928
rect 6135 8925 6147 8959
rect 6089 8919 6147 8925
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6880 8928 7297 8956
rect 6880 8916 6886 8928
rect 7285 8925 7297 8928
rect 7331 8925 7343 8959
rect 7285 8919 7343 8925
rect 8110 8916 8116 8968
rect 8168 8956 8174 8968
rect 8205 8959 8263 8965
rect 8205 8956 8217 8959
rect 8168 8928 8217 8956
rect 8168 8916 8174 8928
rect 8205 8925 8217 8928
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8386 8916 8392 8968
rect 8444 8916 8450 8968
rect 5337 8891 5396 8897
rect 5337 8888 5349 8891
rect 4856 8860 5349 8888
rect 4856 8848 4862 8860
rect 5337 8857 5349 8860
rect 5383 8860 5396 8891
rect 5383 8857 5395 8860
rect 5337 8851 5395 8857
rect 5534 8848 5540 8900
rect 5592 8848 5598 8900
rect 5994 8848 6000 8900
rect 6052 8848 6058 8900
rect 6380 8888 6408 8916
rect 6730 8888 6736 8900
rect 6104 8860 6316 8888
rect 6380 8860 6736 8888
rect 3988 8792 4384 8820
rect 3329 8783 3387 8789
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4706 8820 4712 8832
rect 4488 8792 4712 8820
rect 4488 8780 4494 8792
rect 4706 8780 4712 8792
rect 4764 8820 4770 8832
rect 5810 8829 5816 8832
rect 5629 8823 5687 8829
rect 5629 8820 5641 8823
rect 4764 8792 5641 8820
rect 4764 8780 4770 8792
rect 5629 8789 5641 8792
rect 5675 8789 5687 8823
rect 5629 8783 5687 8789
rect 5792 8823 5816 8829
rect 5792 8789 5804 8823
rect 5868 8820 5874 8832
rect 6104 8820 6132 8860
rect 5868 8792 6132 8820
rect 5792 8783 5816 8789
rect 5810 8780 5816 8783
rect 5868 8780 5874 8792
rect 6178 8780 6184 8832
rect 6236 8780 6242 8832
rect 6288 8820 6316 8860
rect 6730 8848 6736 8860
rect 6788 8848 6794 8900
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7653 8891 7711 8897
rect 7653 8888 7665 8891
rect 7248 8860 7665 8888
rect 7248 8848 7254 8860
rect 7653 8857 7665 8860
rect 7699 8857 7711 8891
rect 7653 8851 7711 8857
rect 9214 8848 9220 8900
rect 9272 8888 9278 8900
rect 9309 8891 9367 8897
rect 9309 8888 9321 8891
rect 9272 8860 9321 8888
rect 9272 8848 9278 8860
rect 9309 8857 9321 8860
rect 9355 8857 9367 8891
rect 9309 8851 9367 8857
rect 10318 8848 10324 8900
rect 10376 8848 10382 8900
rect 6546 8820 6552 8832
rect 6288 8792 6552 8820
rect 6546 8780 6552 8792
rect 6604 8780 6610 8832
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 9122 8780 9128 8832
rect 9180 8820 9186 8832
rect 9674 8820 9680 8832
rect 9180 8792 9680 8820
rect 9180 8780 9186 8792
rect 9674 8780 9680 8792
rect 9732 8780 9738 8832
rect 9950 8780 9956 8832
rect 10008 8820 10014 8832
rect 10781 8823 10839 8829
rect 10781 8820 10793 8823
rect 10008 8792 10793 8820
rect 10008 8780 10014 8792
rect 10781 8789 10793 8792
rect 10827 8789 10839 8823
rect 10781 8783 10839 8789
rect 1104 8730 11224 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 11224 8730
rect 1104 8656 11224 8678
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8616 5043 8619
rect 5442 8616 5448 8628
rect 5031 8588 5448 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5534 8576 5540 8628
rect 5592 8616 5598 8628
rect 6086 8616 6092 8628
rect 5592 8588 6092 8616
rect 5592 8576 5598 8588
rect 6086 8576 6092 8588
rect 6144 8576 6150 8628
rect 8938 8616 8944 8628
rect 6840 8588 8944 8616
rect 4617 8551 4675 8557
rect 4617 8517 4629 8551
rect 4663 8548 4675 8551
rect 6638 8548 6644 8560
rect 4663 8520 6644 8548
rect 4663 8517 4675 8520
rect 4617 8511 4675 8517
rect 6638 8508 6644 8520
rect 6696 8508 6702 8560
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 3142 8480 3148 8492
rect 1719 8452 3148 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 4522 8440 4528 8492
rect 4580 8480 4586 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4580 8452 4905 8480
rect 4580 8440 4586 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 4893 8443 4951 8449
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5353 8483 5411 8489
rect 5215 8452 5304 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 1394 8372 1400 8424
rect 1452 8412 1458 8424
rect 2038 8412 2044 8424
rect 1452 8384 2044 8412
rect 1452 8372 1458 8384
rect 2038 8372 2044 8384
rect 2096 8412 2102 8424
rect 2869 8415 2927 8421
rect 2869 8412 2881 8415
rect 2096 8384 2881 8412
rect 2096 8372 2102 8384
rect 2869 8381 2881 8384
rect 2915 8381 2927 8415
rect 2869 8375 2927 8381
rect 1486 8304 1492 8356
rect 1544 8304 1550 8356
rect 4614 8304 4620 8356
rect 4672 8344 4678 8356
rect 4801 8347 4859 8353
rect 4801 8344 4813 8347
rect 4672 8316 4813 8344
rect 4672 8304 4678 8316
rect 4801 8313 4813 8316
rect 4847 8313 4859 8347
rect 4908 8344 4936 8443
rect 5276 8344 5304 8452
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5810 8480 5816 8492
rect 5399 8452 5816 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6089 8483 6147 8489
rect 6089 8449 6101 8483
rect 6135 8449 6147 8483
rect 6089 8443 6147 8449
rect 5442 8372 5448 8424
rect 5500 8412 5506 8424
rect 5537 8415 5595 8421
rect 5537 8412 5549 8415
rect 5500 8384 5549 8412
rect 5500 8372 5506 8384
rect 5537 8381 5549 8384
rect 5583 8381 5595 8415
rect 5537 8375 5595 8381
rect 5626 8372 5632 8424
rect 5684 8412 5690 8424
rect 6104 8412 6132 8443
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6840 8489 6868 8588
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9033 8619 9091 8625
rect 9033 8585 9045 8619
rect 9079 8616 9091 8619
rect 9122 8616 9128 8628
rect 9079 8588 9128 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9364 8588 9628 8616
rect 9364 8576 9370 8588
rect 7834 8508 7840 8560
rect 7892 8508 7898 8560
rect 9600 8499 9628 8588
rect 9674 8576 9680 8628
rect 9732 8576 9738 8628
rect 10318 8576 10324 8628
rect 10376 8576 10382 8628
rect 9585 8493 9643 8499
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6328 8452 6377 8480
rect 6328 8440 6334 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 6825 8443 6883 8449
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9306 8480 9312 8492
rect 8904 8452 9312 8480
rect 8904 8440 8910 8452
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 9398 8440 9404 8492
rect 9456 8480 9462 8492
rect 9493 8483 9551 8489
rect 9493 8480 9505 8483
rect 9456 8452 9505 8480
rect 9456 8440 9462 8452
rect 9493 8449 9505 8452
rect 9539 8449 9551 8483
rect 9585 8459 9597 8493
rect 9631 8459 9643 8493
rect 9585 8453 9643 8459
rect 9769 8483 9827 8489
rect 9493 8443 9551 8449
rect 9769 8449 9781 8483
rect 9815 8480 9827 8483
rect 9950 8480 9956 8492
rect 9815 8452 9956 8480
rect 9815 8449 9827 8452
rect 9769 8443 9827 8449
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 10226 8440 10232 8492
rect 10284 8440 10290 8492
rect 5684 8384 6868 8412
rect 5684 8372 5690 8384
rect 6840 8356 6868 8384
rect 7098 8372 7104 8424
rect 7156 8372 7162 8424
rect 8110 8372 8116 8424
rect 8168 8412 8174 8424
rect 8864 8412 8892 8440
rect 8168 8384 8892 8412
rect 8168 8372 8174 8384
rect 6730 8344 6736 8356
rect 4908 8316 5212 8344
rect 5276 8316 6736 8344
rect 4801 8307 4859 8313
rect 5184 8276 5212 8316
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 6822 8304 6828 8356
rect 6880 8304 6886 8356
rect 8570 8304 8576 8356
rect 8628 8304 8634 8356
rect 8665 8347 8723 8353
rect 8665 8313 8677 8347
rect 8711 8344 8723 8347
rect 9309 8347 9367 8353
rect 9309 8344 9321 8347
rect 8711 8316 9321 8344
rect 8711 8313 8723 8316
rect 8665 8307 8723 8313
rect 9309 8313 9321 8316
rect 9355 8313 9367 8347
rect 9309 8307 9367 8313
rect 9628 8304 9634 8356
rect 9686 8344 9692 8356
rect 10042 8344 10048 8356
rect 9686 8316 10048 8344
rect 9686 8304 9692 8316
rect 10042 8304 10048 8316
rect 10100 8304 10106 8356
rect 5718 8276 5724 8288
rect 5184 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8276 5782 8288
rect 6270 8276 6276 8288
rect 5776 8248 6276 8276
rect 5776 8236 5782 8248
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 6457 8279 6515 8285
rect 6457 8276 6469 8279
rect 6420 8248 6469 8276
rect 6420 8236 6426 8248
rect 6457 8245 6469 8248
rect 6503 8245 6515 8279
rect 6457 8239 6515 8245
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 9033 8279 9091 8285
rect 9033 8276 9045 8279
rect 7248 8248 9045 8276
rect 7248 8236 7254 8248
rect 9033 8245 9045 8248
rect 9079 8276 9091 8279
rect 9214 8276 9220 8288
rect 9079 8248 9220 8276
rect 9079 8245 9091 8248
rect 9033 8239 9091 8245
rect 9214 8236 9220 8248
rect 9272 8236 9278 8288
rect 1104 8186 11224 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 11224 8186
rect 1104 8112 11224 8134
rect 3142 8032 3148 8084
rect 3200 8032 3206 8084
rect 6730 8032 6736 8084
rect 6788 8032 6794 8084
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 7650 8032 7656 8084
rect 7708 8032 7714 8084
rect 7834 8032 7840 8084
rect 7892 8072 7898 8084
rect 7929 8075 7987 8081
rect 7929 8072 7941 8075
rect 7892 8044 7941 8072
rect 7892 8032 7898 8044
rect 7929 8041 7941 8044
rect 7975 8041 7987 8075
rect 7929 8035 7987 8041
rect 4617 8007 4675 8013
rect 4617 8004 4629 8007
rect 3436 7976 4629 8004
rect 2682 7896 2688 7948
rect 2740 7936 2746 7948
rect 3237 7939 3295 7945
rect 3237 7936 3249 7939
rect 2740 7908 3249 7936
rect 2740 7896 2746 7908
rect 3237 7905 3249 7908
rect 3283 7936 3295 7939
rect 3326 7936 3332 7948
rect 3283 7908 3332 7936
rect 3283 7905 3295 7908
rect 3237 7899 3295 7905
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 3436 7877 3464 7976
rect 4617 7973 4629 7976
rect 4663 7973 4675 8007
rect 4617 7967 4675 7973
rect 6546 7964 6552 8016
rect 6604 8004 6610 8016
rect 6825 8007 6883 8013
rect 6825 8004 6837 8007
rect 6604 7976 6837 8004
rect 6604 7964 6610 7976
rect 6825 7973 6837 7976
rect 6871 7973 6883 8007
rect 6825 7967 6883 7973
rect 7098 7964 7104 8016
rect 7156 8004 7162 8016
rect 7377 8007 7435 8013
rect 7377 8004 7389 8007
rect 7156 7976 7389 8004
rect 7156 7964 7162 7976
rect 7377 7973 7389 7976
rect 7423 7973 7435 8007
rect 7377 7967 7435 7973
rect 3510 7896 3516 7948
rect 3568 7936 3574 7948
rect 3881 7939 3939 7945
rect 3881 7936 3893 7939
rect 3568 7908 3893 7936
rect 3568 7896 3574 7908
rect 3881 7905 3893 7908
rect 3927 7905 3939 7939
rect 3881 7899 3939 7905
rect 4154 7896 4160 7948
rect 4212 7936 4218 7948
rect 4985 7939 5043 7945
rect 4985 7936 4997 7939
rect 4212 7908 4997 7936
rect 4212 7896 4218 7908
rect 4985 7905 4997 7908
rect 5031 7905 5043 7939
rect 4985 7899 5043 7905
rect 5258 7896 5264 7948
rect 5316 7896 5322 7948
rect 8294 7936 8300 7948
rect 7760 7908 8300 7936
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 4433 7871 4491 7877
rect 4433 7837 4445 7871
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 4617 7871 4675 7877
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4706 7868 4712 7880
rect 4663 7840 4712 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 1578 7760 1584 7812
rect 1636 7800 1642 7812
rect 1673 7803 1731 7809
rect 1673 7800 1685 7803
rect 1636 7772 1685 7800
rect 1636 7760 1642 7772
rect 1673 7769 1685 7772
rect 1719 7769 1731 7803
rect 3326 7800 3332 7812
rect 2898 7772 3332 7800
rect 1673 7763 1731 7769
rect 3326 7760 3332 7772
rect 3384 7760 3390 7812
rect 4448 7800 4476 7831
rect 4706 7828 4712 7840
rect 4764 7828 4770 7880
rect 4798 7828 4804 7880
rect 4856 7868 4862 7880
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4856 7840 4905 7868
rect 4856 7828 4862 7840
rect 4893 7837 4905 7840
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 7760 7877 7788 7908
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 7745 7831 7803 7837
rect 7834 7828 7840 7880
rect 7892 7828 7898 7880
rect 5534 7800 5540 7812
rect 4448 7772 5540 7800
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 7193 7803 7251 7809
rect 7193 7769 7205 7803
rect 7239 7800 7251 7803
rect 8018 7800 8024 7812
rect 7239 7772 8024 7800
rect 7239 7769 7251 7772
rect 7193 7763 7251 7769
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 3510 7692 3516 7744
rect 3568 7732 3574 7744
rect 3605 7735 3663 7741
rect 3605 7732 3617 7735
rect 3568 7704 3617 7732
rect 3568 7692 3574 7704
rect 3605 7701 3617 7704
rect 3651 7701 3663 7735
rect 3605 7695 3663 7701
rect 4801 7735 4859 7741
rect 4801 7701 4813 7735
rect 4847 7732 4859 7735
rect 6178 7732 6184 7744
rect 4847 7704 6184 7732
rect 4847 7701 4859 7704
rect 4801 7695 4859 7701
rect 6178 7692 6184 7704
rect 6236 7692 6242 7744
rect 1104 7642 11224 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 11224 7642
rect 1104 7568 11224 7590
rect 3326 7488 3332 7540
rect 3384 7488 3390 7540
rect 5353 7531 5411 7537
rect 5353 7497 5365 7531
rect 5399 7528 5411 7531
rect 5994 7528 6000 7540
rect 5399 7500 6000 7528
rect 5399 7497 5411 7500
rect 5353 7491 5411 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 9030 7488 9036 7540
rect 9088 7528 9094 7540
rect 9309 7531 9367 7537
rect 9309 7528 9321 7531
rect 9088 7500 9321 7528
rect 9088 7488 9094 7500
rect 9309 7497 9321 7500
rect 9355 7497 9367 7531
rect 9309 7491 9367 7497
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 4154 7460 4160 7472
rect 1544 7432 4160 7460
rect 1544 7420 1550 7432
rect 1765 7395 1823 7401
rect 1765 7361 1777 7395
rect 1811 7392 1823 7395
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 1811 7364 2513 7392
rect 1811 7361 1823 7364
rect 1765 7355 1823 7361
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 3142 7352 3148 7404
rect 3200 7352 3206 7404
rect 3620 7401 3648 7432
rect 4154 7420 4160 7432
rect 4212 7420 4218 7472
rect 4614 7420 4620 7472
rect 4672 7420 4678 7472
rect 6638 7420 6644 7472
rect 6696 7460 6702 7472
rect 8021 7463 8079 7469
rect 8021 7460 8033 7463
rect 6696 7432 8033 7460
rect 6696 7420 6702 7432
rect 8021 7429 8033 7432
rect 8067 7429 8079 7463
rect 8021 7423 8079 7429
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 3605 7395 3663 7401
rect 3605 7361 3617 7395
rect 3651 7361 3663 7395
rect 3605 7355 3663 7361
rect 1857 7327 1915 7333
rect 1857 7293 1869 7327
rect 1903 7324 1915 7327
rect 2682 7324 2688 7336
rect 1903 7296 2688 7324
rect 1903 7293 1915 7296
rect 1857 7287 1915 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 1397 7259 1455 7265
rect 1397 7225 1409 7259
rect 1443 7256 1455 7259
rect 1578 7256 1584 7268
rect 1443 7228 1584 7256
rect 1443 7225 1455 7228
rect 1397 7219 1455 7225
rect 1578 7216 1584 7228
rect 1636 7216 1642 7268
rect 3436 7256 3464 7355
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 9030 7392 9036 7404
rect 7883 7364 9036 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 9030 7352 9036 7364
rect 9088 7352 9094 7404
rect 3510 7284 3516 7336
rect 3568 7324 3574 7336
rect 3881 7327 3939 7333
rect 3881 7324 3893 7327
rect 3568 7296 3893 7324
rect 3568 7284 3574 7296
rect 3881 7293 3893 7296
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 3602 7256 3608 7268
rect 3436 7228 3608 7256
rect 3602 7216 3608 7228
rect 3660 7216 3666 7268
rect 5810 7148 5816 7200
rect 5868 7148 5874 7200
rect 1104 7098 11224 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 11224 7098
rect 1104 7024 11224 7046
rect 6638 6944 6644 6996
rect 6696 6944 6702 6996
rect 7190 6944 7196 6996
rect 7248 6984 7254 6996
rect 7377 6987 7435 6993
rect 7377 6984 7389 6987
rect 7248 6956 7389 6984
rect 7248 6944 7254 6956
rect 7377 6953 7389 6956
rect 7423 6953 7435 6987
rect 7377 6947 7435 6953
rect 8864 6888 9076 6916
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 1765 6851 1823 6857
rect 1765 6848 1777 6851
rect 1544 6820 1777 6848
rect 1544 6808 1550 6820
rect 1765 6817 1777 6820
rect 1811 6817 1823 6851
rect 1765 6811 1823 6817
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 3973 6783 4031 6789
rect 3973 6780 3985 6783
rect 3752 6752 3985 6780
rect 3752 6740 3758 6752
rect 3973 6749 3985 6752
rect 4019 6749 4031 6783
rect 3973 6743 4031 6749
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 7742 6740 7748 6792
rect 7800 6740 7806 6792
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 7892 6752 8033 6780
rect 7892 6740 7898 6752
rect 8021 6749 8033 6752
rect 8067 6780 8079 6783
rect 8864 6780 8892 6888
rect 8938 6808 8944 6860
rect 8996 6808 9002 6860
rect 9048 6848 9076 6888
rect 10226 6848 10232 6860
rect 9048 6820 10232 6848
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 8067 6752 8892 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 2038 6672 2044 6724
rect 2096 6672 2102 6724
rect 3881 6715 3939 6721
rect 3881 6712 3893 6715
rect 3266 6684 3893 6712
rect 3881 6681 3893 6684
rect 3927 6681 3939 6715
rect 3881 6675 3939 6681
rect 9214 6672 9220 6724
rect 9272 6672 9278 6724
rect 10226 6672 10232 6724
rect 10284 6672 10290 6724
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 3513 6647 3571 6653
rect 3513 6644 3525 6647
rect 2924 6616 3525 6644
rect 2924 6604 2930 6616
rect 3513 6613 3525 6616
rect 3559 6613 3571 6647
rect 3513 6607 3571 6613
rect 7190 6604 7196 6656
rect 7248 6604 7254 6656
rect 7374 6604 7380 6656
rect 7432 6604 7438 6656
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7524 6616 7941 6644
rect 7524 6604 7530 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 9548 6616 10701 6644
rect 9548 6604 9554 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 1104 6554 11224 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 11224 6554
rect 1104 6480 11224 6502
rect 2038 6400 2044 6452
rect 2096 6440 2102 6452
rect 2133 6443 2191 6449
rect 2133 6440 2145 6443
rect 2096 6412 2145 6440
rect 2096 6400 2102 6412
rect 2133 6409 2145 6412
rect 2179 6409 2191 6443
rect 2133 6403 2191 6409
rect 7190 6400 7196 6452
rect 7248 6440 7254 6452
rect 7248 6412 7972 6440
rect 7248 6400 7254 6412
rect 2593 6375 2651 6381
rect 2593 6341 2605 6375
rect 2639 6372 2651 6375
rect 2866 6372 2872 6384
rect 2639 6344 2872 6372
rect 2639 6341 2651 6344
rect 2593 6335 2651 6341
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 4614 6332 4620 6384
rect 4672 6372 4678 6384
rect 5873 6375 5931 6381
rect 5873 6372 5885 6375
rect 4672 6344 5885 6372
rect 4672 6332 4678 6344
rect 5873 6341 5885 6344
rect 5919 6341 5931 6375
rect 5873 6335 5931 6341
rect 6086 6332 6092 6384
rect 6144 6332 6150 6384
rect 7466 6332 7472 6384
rect 7524 6332 7530 6384
rect 7944 6381 7972 6412
rect 8018 6400 8024 6452
rect 8076 6440 8082 6452
rect 8481 6443 8539 6449
rect 8481 6440 8493 6443
rect 8076 6412 8493 6440
rect 8076 6400 8082 6412
rect 8481 6409 8493 6412
rect 8527 6409 8539 6443
rect 8481 6403 8539 6409
rect 8846 6400 8852 6452
rect 8904 6400 8910 6452
rect 9214 6400 9220 6452
rect 9272 6440 9278 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 9272 6412 9505 6440
rect 9272 6400 9278 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 10137 6443 10195 6449
rect 10137 6409 10149 6443
rect 10183 6440 10195 6443
rect 10226 6440 10232 6452
rect 10183 6412 10232 6440
rect 10183 6409 10195 6412
rect 10137 6403 10195 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 7929 6375 7987 6381
rect 7929 6341 7941 6375
rect 7975 6341 7987 6375
rect 8938 6372 8944 6384
rect 7929 6335 7987 6341
rect 8220 6344 8944 6372
rect 1486 6264 1492 6316
rect 1544 6304 1550 6316
rect 2685 6307 2743 6313
rect 2685 6304 2697 6307
rect 1544 6276 2697 6304
rect 1544 6264 1550 6276
rect 2685 6273 2697 6276
rect 2731 6273 2743 6307
rect 2685 6267 2743 6273
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5261 6307 5319 6313
rect 5261 6304 5273 6307
rect 5224 6276 5273 6304
rect 5224 6264 5230 6276
rect 5261 6273 5273 6276
rect 5307 6273 5319 6307
rect 5261 6267 5319 6273
rect 5445 6307 5503 6313
rect 5445 6273 5457 6307
rect 5491 6304 5503 6307
rect 6454 6304 6460 6316
rect 5491 6276 6460 6304
rect 5491 6273 5503 6276
rect 5445 6267 5503 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 8220 6313 8248 6344
rect 8938 6332 8944 6344
rect 8996 6332 9002 6384
rect 9309 6375 9367 6381
rect 9309 6341 9321 6375
rect 9355 6372 9367 6375
rect 9953 6375 10011 6381
rect 9953 6372 9965 6375
rect 9355 6344 9965 6372
rect 9355 6341 9367 6344
rect 9309 6335 9367 6341
rect 9953 6341 9965 6344
rect 9999 6341 10011 6375
rect 9953 6335 10011 6341
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6273 8263 6307
rect 8205 6267 8263 6273
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8570 6264 8576 6316
rect 8628 6264 8634 6316
rect 8662 6264 8668 6316
rect 8720 6264 8726 6316
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 9585 6307 9643 6313
rect 9585 6304 9597 6307
rect 8812 6276 9597 6304
rect 8812 6264 8818 6276
rect 9585 6273 9597 6276
rect 9631 6273 9643 6307
rect 9585 6267 9643 6273
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10229 6307 10287 6313
rect 10229 6273 10241 6307
rect 10275 6304 10287 6307
rect 10318 6304 10324 6316
rect 10275 6276 10324 6304
rect 10275 6273 10287 6276
rect 10229 6267 10287 6273
rect 2961 6239 3019 6245
rect 2961 6205 2973 6239
rect 3007 6236 3019 6239
rect 3050 6236 3056 6248
rect 3007 6208 3056 6236
rect 3007 6205 3019 6208
rect 2961 6199 3019 6205
rect 3050 6196 3056 6208
rect 3108 6196 3114 6248
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 5350 6236 5356 6248
rect 3660 6208 5356 6236
rect 3660 6196 3666 6208
rect 5350 6196 5356 6208
rect 5408 6236 5414 6248
rect 6086 6236 6092 6248
rect 5408 6208 6092 6236
rect 5408 6196 5414 6208
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 8312 6236 8340 6264
rect 9490 6236 9496 6248
rect 8312 6208 9496 6236
rect 9490 6196 9496 6208
rect 9548 6236 9554 6248
rect 9784 6236 9812 6267
rect 10318 6264 10324 6276
rect 10376 6264 10382 6316
rect 9548 6208 9812 6236
rect 9548 6196 9554 6208
rect 2317 6171 2375 6177
rect 2317 6137 2329 6171
rect 2363 6137 2375 6171
rect 2317 6131 2375 6137
rect 5629 6171 5687 6177
rect 5629 6137 5641 6171
rect 5675 6168 5687 6171
rect 5675 6140 5948 6168
rect 5675 6137 5687 6140
rect 5629 6131 5687 6137
rect 2332 6100 2360 6131
rect 3602 6100 3608 6112
rect 2332 6072 3608 6100
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 3694 6060 3700 6112
rect 3752 6100 3758 6112
rect 4433 6103 4491 6109
rect 4433 6100 4445 6103
rect 3752 6072 4445 6100
rect 3752 6060 3758 6072
rect 4433 6069 4445 6072
rect 4479 6100 4491 6103
rect 4706 6100 4712 6112
rect 4479 6072 4712 6100
rect 4479 6069 4491 6072
rect 4433 6063 4491 6069
rect 4706 6060 4712 6072
rect 4764 6060 4770 6112
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 5920 6109 5948 6140
rect 8846 6128 8852 6180
rect 8904 6168 8910 6180
rect 8941 6171 8999 6177
rect 8941 6168 8953 6171
rect 8904 6140 8953 6168
rect 8904 6128 8910 6140
rect 8941 6137 8953 6140
rect 8987 6137 8999 6171
rect 8941 6131 8999 6137
rect 5721 6103 5779 6109
rect 5721 6100 5733 6103
rect 5132 6072 5733 6100
rect 5132 6060 5138 6072
rect 5721 6069 5733 6072
rect 5767 6069 5779 6103
rect 5721 6063 5779 6069
rect 5905 6103 5963 6109
rect 5905 6069 5917 6103
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 6914 6100 6920 6112
rect 6503 6072 6920 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 9306 6060 9312 6112
rect 9364 6060 9370 6112
rect 1104 6010 11224 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 11224 6010
rect 1104 5936 11224 5958
rect 3050 5856 3056 5908
rect 3108 5856 3114 5908
rect 3237 5899 3295 5905
rect 3237 5865 3249 5899
rect 3283 5865 3295 5899
rect 3237 5859 3295 5865
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 3970 5896 3976 5908
rect 3927 5868 3976 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 2961 5831 3019 5837
rect 2961 5797 2973 5831
rect 3007 5828 3019 5831
rect 3252 5828 3280 5859
rect 3970 5856 3976 5868
rect 4028 5856 4034 5908
rect 4614 5856 4620 5908
rect 4672 5856 4678 5908
rect 5166 5896 5172 5908
rect 4724 5868 5172 5896
rect 4724 5828 4752 5868
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 7193 5899 7251 5905
rect 7193 5865 7205 5899
rect 7239 5896 7251 5899
rect 7374 5896 7380 5908
rect 7239 5868 7380 5896
rect 7239 5865 7251 5868
rect 7193 5859 7251 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7653 5899 7711 5905
rect 7653 5865 7665 5899
rect 7699 5896 7711 5899
rect 7742 5896 7748 5908
rect 7699 5868 7748 5896
rect 7699 5865 7711 5868
rect 7653 5859 7711 5865
rect 7742 5856 7748 5868
rect 7800 5856 7806 5908
rect 8113 5899 8171 5905
rect 8113 5865 8125 5899
rect 8159 5896 8171 5899
rect 8570 5896 8576 5908
rect 8159 5868 8576 5896
rect 8159 5865 8171 5868
rect 8113 5859 8171 5865
rect 8018 5828 8024 5840
rect 3007 5800 3280 5828
rect 4540 5800 4752 5828
rect 7300 5800 8024 5828
rect 3007 5797 3019 5800
rect 2961 5791 3019 5797
rect 2866 5760 2872 5772
rect 2332 5732 2872 5760
rect 2332 5701 2360 5732
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2501 5695 2559 5701
rect 2501 5661 2513 5695
rect 2547 5692 2559 5695
rect 2682 5692 2688 5704
rect 2547 5664 2688 5692
rect 2547 5661 2559 5664
rect 2501 5655 2559 5661
rect 2332 5624 2360 5655
rect 2682 5652 2688 5664
rect 2740 5692 2746 5704
rect 2777 5695 2835 5701
rect 2777 5692 2789 5695
rect 2740 5664 2789 5692
rect 2740 5652 2746 5664
rect 2777 5661 2789 5664
rect 2823 5692 2835 5695
rect 3694 5692 3700 5704
rect 2823 5664 3700 5692
rect 2823 5661 2835 5664
rect 2777 5655 2835 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3844 5664 3985 5692
rect 3844 5652 3850 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4246 5652 4252 5704
rect 4304 5692 4310 5704
rect 4540 5701 4568 5800
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 4801 5763 4859 5769
rect 4801 5760 4813 5763
rect 4672 5732 4813 5760
rect 4672 5720 4678 5732
rect 4801 5729 4813 5732
rect 4847 5729 4859 5763
rect 4801 5723 4859 5729
rect 5074 5720 5080 5772
rect 5132 5720 5138 5772
rect 5166 5720 5172 5772
rect 5224 5760 5230 5772
rect 7300 5769 7328 5800
rect 8018 5788 8024 5800
rect 8076 5788 8082 5840
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 5224 5732 7297 5760
rect 5224 5720 5230 5732
rect 6748 5701 6776 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 8128 5760 8156 5859
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 8665 5899 8723 5905
rect 8665 5865 8677 5899
rect 8711 5896 8723 5899
rect 8754 5896 8760 5908
rect 8711 5868 8760 5896
rect 8711 5865 8723 5868
rect 8665 5859 8723 5865
rect 8478 5788 8484 5840
rect 8536 5828 8542 5840
rect 8680 5828 8708 5859
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5865 9183 5899
rect 9125 5859 9183 5865
rect 8536 5800 8708 5828
rect 8536 5788 8542 5800
rect 7285 5723 7343 5729
rect 7484 5732 8156 5760
rect 4525 5695 4583 5701
rect 4525 5692 4537 5695
rect 4304 5664 4537 5692
rect 4304 5652 4310 5664
rect 4525 5661 4537 5664
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4709 5695 4767 5701
rect 4709 5661 4721 5695
rect 4755 5661 4767 5695
rect 4709 5655 4767 5661
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5661 6791 5695
rect 6733 5655 6791 5661
rect 2593 5627 2651 5633
rect 2593 5624 2605 5627
rect 2332 5596 2605 5624
rect 2593 5593 2605 5596
rect 2639 5593 2651 5627
rect 3205 5627 3263 5633
rect 3205 5624 3217 5627
rect 2593 5587 2651 5593
rect 2884 5596 3217 5624
rect 2501 5559 2559 5565
rect 2501 5525 2513 5559
rect 2547 5556 2559 5559
rect 2884 5556 2912 5596
rect 3205 5593 3217 5596
rect 3251 5593 3263 5627
rect 3205 5587 3263 5593
rect 3418 5584 3424 5636
rect 3476 5584 3482 5636
rect 2547 5528 2912 5556
rect 4724 5556 4752 5655
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6972 5664 7021 5692
rect 6972 5652 6978 5664
rect 7009 5661 7021 5664
rect 7055 5692 7067 5695
rect 7098 5692 7104 5704
rect 7055 5664 7104 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7484 5701 7512 5732
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5661 7803 5695
rect 7745 5655 7803 5661
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5692 8539 5695
rect 8570 5692 8576 5704
rect 8527 5664 8576 5692
rect 8527 5661 8539 5664
rect 8481 5655 8539 5661
rect 5810 5584 5816 5636
rect 5868 5584 5874 5636
rect 7116 5624 7144 5652
rect 7760 5624 7788 5655
rect 7116 5596 7788 5624
rect 6454 5556 6460 5568
rect 4724 5528 6460 5556
rect 2547 5525 2559 5528
rect 2501 5519 2559 5525
rect 6454 5516 6460 5528
rect 6512 5556 6518 5568
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 6512 5528 6561 5556
rect 6512 5516 6518 5528
rect 6549 5525 6561 5528
rect 6595 5556 6607 5559
rect 6825 5559 6883 5565
rect 6825 5556 6837 5559
rect 6595 5528 6837 5556
rect 6595 5525 6607 5528
rect 6549 5519 6607 5525
rect 6825 5525 6837 5528
rect 6871 5556 6883 5559
rect 7944 5556 7972 5655
rect 8570 5652 8576 5664
rect 8628 5652 8634 5704
rect 8665 5695 8723 5701
rect 8665 5661 8677 5695
rect 8711 5692 8723 5695
rect 9140 5692 9168 5859
rect 10318 5856 10324 5908
rect 10376 5856 10382 5908
rect 8711 5664 9168 5692
rect 8711 5661 8723 5664
rect 8665 5655 8723 5661
rect 8294 5584 8300 5636
rect 8352 5624 8358 5636
rect 8680 5624 8708 5655
rect 9306 5652 9312 5704
rect 9364 5652 9370 5704
rect 9953 5695 10011 5701
rect 9953 5661 9965 5695
rect 9999 5692 10011 5695
rect 10318 5692 10324 5704
rect 9999 5664 10324 5692
rect 9999 5661 10011 5664
rect 9953 5655 10011 5661
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 8352 5596 8708 5624
rect 8941 5627 8999 5633
rect 8352 5584 8358 5596
rect 8941 5593 8953 5627
rect 8987 5624 8999 5627
rect 9030 5624 9036 5636
rect 8987 5596 9036 5624
rect 8987 5593 8999 5596
rect 8941 5587 8999 5593
rect 9030 5584 9036 5596
rect 9088 5624 9094 5636
rect 9324 5624 9352 5652
rect 9088 5596 9352 5624
rect 9088 5584 9094 5596
rect 10410 5584 10416 5636
rect 10468 5624 10474 5636
rect 10597 5627 10655 5633
rect 10597 5624 10609 5627
rect 10468 5596 10609 5624
rect 10468 5584 10474 5596
rect 10597 5593 10609 5596
rect 10643 5593 10655 5627
rect 10597 5587 10655 5593
rect 6871 5528 7972 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 9141 5559 9199 5565
rect 9141 5556 9153 5559
rect 8812 5528 9153 5556
rect 8812 5516 8818 5528
rect 9141 5525 9153 5528
rect 9187 5525 9199 5559
rect 9141 5519 9199 5525
rect 9306 5516 9312 5568
rect 9364 5516 9370 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 1104 5466 11224 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 11224 5466
rect 1104 5392 11224 5414
rect 2301 5355 2359 5361
rect 2301 5321 2313 5355
rect 2347 5352 2359 5355
rect 2593 5355 2651 5361
rect 2593 5352 2605 5355
rect 2347 5324 2605 5352
rect 2347 5321 2359 5324
rect 2301 5315 2359 5321
rect 2593 5321 2605 5324
rect 2639 5321 2651 5355
rect 2593 5315 2651 5321
rect 4246 5312 4252 5364
rect 4304 5312 4310 5364
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 4706 5352 4712 5364
rect 4571 5324 4712 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8294 5352 8300 5364
rect 7975 5324 8300 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 8389 5355 8447 5361
rect 8389 5321 8401 5355
rect 8435 5352 8447 5355
rect 8662 5352 8668 5364
rect 8435 5324 8668 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 10410 5352 10416 5364
rect 8772 5324 10416 5352
rect 2501 5287 2559 5293
rect 2501 5253 2513 5287
rect 2547 5284 2559 5287
rect 3418 5284 3424 5296
rect 2547 5256 3424 5284
rect 2547 5253 2559 5256
rect 2501 5247 2559 5253
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 3786 5244 3792 5296
rect 3844 5284 3850 5296
rect 5537 5287 5595 5293
rect 5537 5284 5549 5287
rect 3844 5256 5549 5284
rect 3844 5244 3850 5256
rect 5537 5253 5549 5256
rect 5583 5284 5595 5287
rect 5626 5284 5632 5296
rect 5583 5256 5632 5284
rect 5583 5253 5595 5256
rect 5537 5247 5595 5253
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 8772 5284 8800 5324
rect 10410 5312 10416 5324
rect 10468 5312 10474 5364
rect 5828 5256 8800 5284
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 2498 5108 2504 5160
rect 2556 5148 2562 5160
rect 2608 5148 2636 5179
rect 2682 5176 2688 5228
rect 2740 5176 2746 5228
rect 2866 5176 2872 5228
rect 2924 5216 2930 5228
rect 3970 5216 3976 5228
rect 2924 5188 3976 5216
rect 2924 5176 2930 5188
rect 3970 5176 3976 5188
rect 4028 5216 4034 5228
rect 5828 5225 5856 5256
rect 8846 5244 8852 5296
rect 8904 5244 8910 5296
rect 10042 5244 10048 5296
rect 10100 5244 10106 5296
rect 4433 5219 4491 5225
rect 4433 5216 4445 5219
rect 4028 5188 4445 5216
rect 4028 5176 4034 5188
rect 4433 5185 4445 5188
rect 4479 5185 4491 5219
rect 4433 5179 4491 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 4632 5148 4660 5179
rect 7742 5176 7748 5228
rect 7800 5176 7806 5228
rect 7929 5219 7987 5225
rect 7929 5185 7941 5219
rect 7975 5216 7987 5219
rect 8205 5219 8263 5225
rect 8205 5216 8217 5219
rect 7975 5188 8217 5216
rect 7975 5185 7987 5188
rect 7929 5179 7987 5185
rect 8205 5185 8217 5188
rect 8251 5216 8263 5219
rect 8294 5216 8300 5228
rect 8251 5188 8300 5216
rect 8251 5185 8263 5188
rect 8205 5179 8263 5185
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 8478 5176 8484 5228
rect 8536 5176 8542 5228
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9125 5219 9183 5225
rect 9125 5216 9137 5219
rect 8996 5188 9137 5216
rect 8996 5176 9002 5188
rect 9125 5185 9137 5188
rect 9171 5185 9183 5219
rect 9125 5179 9183 5185
rect 2556 5120 4660 5148
rect 8021 5151 8079 5157
rect 2556 5108 2562 5120
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 9401 5151 9459 5157
rect 9401 5148 9413 5151
rect 8067 5120 8984 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 4801 5083 4859 5089
rect 4801 5049 4813 5083
rect 4847 5080 4859 5083
rect 5534 5080 5540 5092
rect 4847 5052 5540 5080
rect 4847 5049 4859 5052
rect 4801 5043 4859 5049
rect 5534 5040 5540 5052
rect 5592 5040 5598 5092
rect 1762 4972 1768 5024
rect 1820 5012 1826 5024
rect 2133 5015 2191 5021
rect 2133 5012 2145 5015
rect 1820 4984 2145 5012
rect 1820 4972 1826 4984
rect 2133 4981 2145 4984
rect 2179 4981 2191 5015
rect 2133 4975 2191 4981
rect 2314 4972 2320 5024
rect 2372 4972 2378 5024
rect 8662 4972 8668 5024
rect 8720 5012 8726 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 8720 4984 8861 5012
rect 8720 4972 8726 4984
rect 8849 4981 8861 4984
rect 8895 4981 8907 5015
rect 8956 5012 8984 5120
rect 9048 5120 9413 5148
rect 9048 5089 9076 5120
rect 9401 5117 9413 5120
rect 9447 5117 9459 5151
rect 9401 5111 9459 5117
rect 9033 5083 9091 5089
rect 9033 5049 9045 5083
rect 9079 5049 9091 5083
rect 9033 5043 9091 5049
rect 9122 5012 9128 5024
rect 8956 4984 9128 5012
rect 8849 4975 8907 4981
rect 9122 4972 9128 4984
rect 9180 5012 9186 5024
rect 10873 5015 10931 5021
rect 10873 5012 10885 5015
rect 9180 4984 10885 5012
rect 9180 4972 9186 4984
rect 10873 4981 10885 4984
rect 10919 4981 10931 5015
rect 10873 4975 10931 4981
rect 1104 4922 11224 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 11224 4922
rect 1104 4848 11224 4870
rect 2498 4768 2504 4820
rect 2556 4808 2562 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 2556 4780 3249 4808
rect 2556 4768 2562 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 8573 4811 8631 4817
rect 8573 4777 8585 4811
rect 8619 4808 8631 4811
rect 8754 4808 8760 4820
rect 8619 4780 8760 4808
rect 8619 4777 8631 4780
rect 8573 4771 8631 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 1486 4632 1492 4684
rect 1544 4672 1550 4684
rect 4341 4675 4399 4681
rect 4341 4672 4353 4675
rect 1544 4644 4353 4672
rect 1544 4632 1550 4644
rect 4341 4641 4353 4644
rect 4387 4672 4399 4675
rect 4614 4672 4620 4684
rect 4387 4644 4620 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 5626 4632 5632 4684
rect 5684 4672 5690 4684
rect 5684 4644 6408 4672
rect 5684 4632 5690 4644
rect 3513 4607 3571 4613
rect 3513 4573 3525 4607
rect 3559 4604 3571 4607
rect 3786 4604 3792 4616
rect 3559 4576 3792 4604
rect 3559 4573 3571 4576
rect 3513 4567 3571 4573
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 6380 4613 6408 4644
rect 8938 4632 8944 4684
rect 8996 4632 9002 4684
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 9306 4672 9312 4684
rect 9263 4644 9312 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 7742 4564 7748 4616
rect 7800 4604 7806 4616
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 7800 4576 8217 4604
rect 7800 4564 7806 4576
rect 8205 4573 8217 4576
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 1762 4496 1768 4548
rect 1820 4496 1826 4548
rect 3421 4539 3479 4545
rect 3421 4536 3433 4539
rect 2990 4508 3433 4536
rect 3421 4505 3433 4508
rect 3467 4505 3479 4539
rect 3421 4499 3479 4505
rect 4617 4539 4675 4545
rect 4617 4505 4629 4539
rect 4663 4536 4675 4539
rect 4706 4536 4712 4548
rect 4663 4508 4712 4536
rect 4663 4505 4675 4508
rect 4617 4499 4675 4505
rect 4706 4496 4712 4508
rect 4764 4496 4770 4548
rect 6273 4539 6331 4545
rect 6273 4536 6285 4539
rect 5842 4508 6285 4536
rect 6273 4505 6285 4508
rect 6319 4505 6331 4539
rect 6273 4499 6331 4505
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4505 8447 4539
rect 8389 4499 8447 4505
rect 5534 4428 5540 4480
rect 5592 4468 5598 4480
rect 5994 4468 6000 4480
rect 5592 4440 6000 4468
rect 5592 4428 5598 4440
rect 5994 4428 6000 4440
rect 6052 4468 6058 4480
rect 6089 4471 6147 4477
rect 6089 4468 6101 4471
rect 6052 4440 6101 4468
rect 6052 4428 6058 4440
rect 6089 4437 6101 4440
rect 6135 4437 6147 4471
rect 6089 4431 6147 4437
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 8404 4468 8432 4499
rect 9950 4496 9956 4548
rect 10008 4496 10014 4548
rect 10689 4471 10747 4477
rect 10689 4468 10701 4471
rect 8352 4440 10701 4468
rect 8352 4428 8358 4440
rect 10689 4437 10701 4440
rect 10735 4437 10747 4471
rect 10689 4431 10747 4437
rect 1104 4378 11224 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 11224 4378
rect 1104 4304 11224 4326
rect 2314 4224 2320 4276
rect 2372 4264 2378 4276
rect 2409 4267 2467 4273
rect 2409 4264 2421 4267
rect 2372 4236 2421 4264
rect 2372 4224 2378 4236
rect 2409 4233 2421 4236
rect 2455 4233 2467 4267
rect 2409 4227 2467 4233
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 2777 4267 2835 4273
rect 2777 4264 2789 4267
rect 2740 4236 2789 4264
rect 2740 4224 2746 4236
rect 2777 4233 2789 4236
rect 2823 4233 2835 4267
rect 2777 4227 2835 4233
rect 4617 4267 4675 4273
rect 4617 4233 4629 4267
rect 4663 4264 4675 4267
rect 4893 4267 4951 4273
rect 4893 4264 4905 4267
rect 4663 4236 4905 4264
rect 4663 4233 4675 4236
rect 4617 4227 4675 4233
rect 4893 4233 4905 4236
rect 4939 4233 4951 4267
rect 4893 4227 4951 4233
rect 8846 4224 8852 4276
rect 8904 4224 8910 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 10468 4236 10701 4264
rect 10468 4224 10474 4236
rect 10689 4233 10701 4236
rect 10735 4233 10747 4267
rect 10689 4227 10747 4233
rect 2608 4168 5304 4196
rect 2498 4088 2504 4140
rect 2556 4128 2562 4140
rect 2608 4137 2636 4168
rect 2593 4131 2651 4137
rect 2593 4128 2605 4131
rect 2556 4100 2605 4128
rect 2556 4088 2562 4100
rect 2593 4097 2605 4100
rect 2639 4097 2651 4131
rect 2593 4091 2651 4097
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 2884 4060 2912 4091
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4249 4131 4307 4137
rect 4249 4128 4261 4131
rect 4212 4100 4261 4128
rect 4212 4088 4218 4100
rect 4249 4097 4261 4100
rect 4295 4097 4307 4131
rect 4249 4091 4307 4097
rect 4798 4088 4804 4140
rect 4856 4128 4862 4140
rect 5276 4137 5304 4168
rect 5534 4156 5540 4208
rect 5592 4156 5598 4208
rect 6825 4199 6883 4205
rect 6825 4165 6837 4199
rect 6871 4196 6883 4199
rect 6871 4168 7236 4196
rect 6871 4165 6883 4168
rect 6825 4159 6883 4165
rect 5169 4131 5227 4137
rect 5169 4128 5181 4131
rect 4856 4100 5181 4128
rect 4856 4088 4862 4100
rect 5169 4097 5181 4100
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 5261 4131 5319 4137
rect 5261 4097 5273 4131
rect 5307 4097 5319 4131
rect 5261 4091 5319 4097
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5552 4128 5580 4156
rect 5399 4100 5580 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 3786 4060 3792 4072
rect 2884 4032 3792 4060
rect 3786 4020 3792 4032
rect 3844 4060 3850 4072
rect 3970 4060 3976 4072
rect 3844 4032 3976 4060
rect 3844 4020 3850 4032
rect 3970 4020 3976 4032
rect 4028 4060 4034 4072
rect 5077 4063 5135 4069
rect 5077 4060 5089 4063
rect 4028 4032 5089 4060
rect 4028 4020 4034 4032
rect 5077 4029 5089 4032
rect 5123 4029 5135 4063
rect 5077 4023 5135 4029
rect 4706 3952 4712 4004
rect 4764 3992 4770 4004
rect 4801 3995 4859 4001
rect 4801 3992 4813 3995
rect 4764 3964 4813 3992
rect 4764 3952 4770 3964
rect 4801 3961 4813 3964
rect 4847 3961 4859 3995
rect 4801 3955 4859 3961
rect 4890 3952 4896 4004
rect 4948 3992 4954 4004
rect 5368 3992 5396 4091
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 7208 4137 7236 4168
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4097 6699 4131
rect 6641 4091 6699 4097
rect 7193 4131 7251 4137
rect 7193 4097 7205 4131
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 6656 4060 6684 4091
rect 7374 4088 7380 4140
rect 7432 4088 7438 4140
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4128 7527 4131
rect 7834 4128 7840 4140
rect 7515 4100 7840 4128
rect 7515 4097 7527 4100
rect 7469 4091 7527 4097
rect 7834 4088 7840 4100
rect 7892 4088 7898 4140
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8444 4100 8677 4128
rect 8444 4088 8450 4100
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8849 4131 8907 4137
rect 8849 4097 8861 4131
rect 8895 4128 8907 4131
rect 9033 4131 9091 4137
rect 9033 4128 9045 4131
rect 8895 4100 9045 4128
rect 8895 4097 8907 4100
rect 8849 4091 8907 4097
rect 9033 4097 9045 4100
rect 9079 4097 9091 4131
rect 9033 4091 9091 4097
rect 5592 4032 6684 4060
rect 7009 4063 7067 4069
rect 5592 4020 5598 4032
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 7558 4060 7564 4072
rect 7055 4032 7564 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 4948 3964 5396 3992
rect 4948 3952 4954 3964
rect 5718 3952 5724 4004
rect 5776 3992 5782 4004
rect 7024 3992 7052 4023
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 8864 4060 8892 4091
rect 9122 4088 9128 4140
rect 9180 4088 9186 4140
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10137 4131 10195 4137
rect 10137 4128 10149 4131
rect 10008 4100 10149 4128
rect 10008 4088 10014 4100
rect 10137 4097 10149 4100
rect 10183 4097 10195 4131
rect 10137 4091 10195 4097
rect 10229 4131 10287 4137
rect 10229 4097 10241 4131
rect 10275 4128 10287 4131
rect 10318 4128 10324 4140
rect 10275 4100 10324 4128
rect 10275 4097 10287 4100
rect 10229 4091 10287 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10870 4088 10876 4140
rect 10928 4088 10934 4140
rect 8628 4032 8892 4060
rect 8628 4020 8634 4032
rect 5776 3964 7052 3992
rect 5776 3952 5782 3964
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 5350 3924 5356 3936
rect 4663 3896 5356 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 6825 3927 6883 3933
rect 6825 3893 6837 3927
rect 6871 3924 6883 3927
rect 7282 3924 7288 3936
rect 6871 3896 7288 3924
rect 6871 3893 6883 3896
rect 6825 3887 6883 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 7984 3896 8217 3924
rect 7984 3884 7990 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8205 3887 8263 3893
rect 1104 3834 11224 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 11224 3834
rect 1104 3760 11224 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 2556 3692 3893 3720
rect 2556 3680 2562 3692
rect 3881 3689 3893 3692
rect 3927 3689 3939 3723
rect 3881 3683 3939 3689
rect 3896 3652 3924 3683
rect 4154 3680 4160 3732
rect 4212 3720 4218 3732
rect 4798 3720 4804 3732
rect 4212 3692 4804 3720
rect 4212 3680 4218 3692
rect 4798 3680 4804 3692
rect 4856 3680 4862 3732
rect 5534 3680 5540 3732
rect 5592 3680 5598 3732
rect 6546 3680 6552 3732
rect 6604 3720 6610 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 6604 3692 6837 3720
rect 6604 3680 6610 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 7374 3680 7380 3732
rect 7432 3720 7438 3732
rect 7653 3723 7711 3729
rect 7653 3720 7665 3723
rect 7432 3692 7665 3720
rect 7432 3680 7438 3692
rect 7653 3689 7665 3692
rect 7699 3689 7711 3723
rect 7653 3683 7711 3689
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3720 8171 3723
rect 8570 3720 8576 3732
rect 8159 3692 8576 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 8570 3680 8576 3692
rect 8628 3680 8634 3732
rect 3896 3624 4292 3652
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 3804 3448 3832 3479
rect 4062 3476 4068 3528
rect 4120 3476 4126 3528
rect 4154 3476 4160 3528
rect 4212 3476 4218 3528
rect 4264 3516 4292 3624
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4387 3556 5028 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4433 3519 4491 3525
rect 4433 3516 4445 3519
rect 4264 3488 4445 3516
rect 4433 3485 4445 3488
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 4890 3516 4896 3528
rect 4847 3488 4896 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5000 3516 5028 3556
rect 5994 3544 6000 3596
rect 6052 3544 6058 3596
rect 5077 3519 5135 3525
rect 5077 3516 5089 3519
rect 5000 3488 5089 3516
rect 5077 3485 5089 3488
rect 5123 3485 5135 3519
rect 5077 3479 5135 3485
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 4522 3448 4528 3460
rect 3804 3420 4528 3448
rect 4522 3408 4528 3420
rect 4580 3448 4586 3460
rect 4617 3451 4675 3457
rect 4617 3448 4629 3451
rect 4580 3420 4629 3448
rect 4580 3408 4586 3420
rect 4617 3417 4629 3420
rect 4663 3417 4675 3451
rect 4617 3411 4675 3417
rect 4706 3408 4712 3460
rect 4764 3408 4770 3460
rect 5368 3448 5396 3479
rect 5718 3476 5724 3528
rect 5776 3476 5782 3528
rect 5902 3476 5908 3528
rect 5960 3476 5966 3528
rect 6086 3476 6092 3528
rect 6144 3476 6150 3528
rect 6273 3519 6331 3525
rect 6273 3485 6285 3519
rect 6319 3516 6331 3519
rect 6546 3516 6552 3528
rect 6319 3488 6552 3516
rect 6319 3485 6331 3488
rect 6273 3479 6331 3485
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 7101 3519 7159 3525
rect 7101 3485 7113 3519
rect 7147 3516 7159 3519
rect 7392 3516 7420 3680
rect 7558 3612 7564 3664
rect 7616 3652 7622 3664
rect 8297 3655 8355 3661
rect 8297 3652 8309 3655
rect 7616 3624 8309 3652
rect 7616 3612 7622 3624
rect 8297 3621 8309 3624
rect 8343 3621 8355 3655
rect 8297 3615 8355 3621
rect 7147 3488 7420 3516
rect 7147 3485 7159 3488
rect 7101 3479 7159 3485
rect 7558 3476 7564 3528
rect 7616 3516 7622 3528
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7616 3488 7849 3516
rect 7616 3476 7622 3488
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3516 8263 3519
rect 8570 3516 8576 3528
rect 8251 3488 8576 3516
rect 8251 3485 8263 3488
rect 8205 3479 8263 3485
rect 8570 3476 8576 3488
rect 8628 3476 8634 3528
rect 8665 3519 8723 3525
rect 8665 3485 8677 3519
rect 8711 3516 8723 3519
rect 9122 3516 9128 3528
rect 8711 3488 9128 3516
rect 8711 3485 8723 3488
rect 8665 3479 8723 3485
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 5000 3420 5396 3448
rect 6457 3451 6515 3457
rect 5000 3389 5028 3420
rect 6457 3417 6469 3451
rect 6503 3448 6515 3451
rect 7377 3451 7435 3457
rect 7377 3448 7389 3451
rect 6503 3420 7389 3448
rect 6503 3417 6515 3420
rect 6457 3411 6515 3417
rect 7377 3417 7389 3420
rect 7423 3417 7435 3451
rect 7377 3411 7435 3417
rect 4985 3383 5043 3389
rect 4985 3349 4997 3383
rect 5031 3349 5043 3383
rect 4985 3343 5043 3349
rect 5169 3383 5227 3389
rect 5169 3349 5181 3383
rect 5215 3380 5227 3383
rect 5258 3380 5264 3392
rect 5215 3352 5264 3380
rect 5215 3349 5227 3352
rect 5169 3343 5227 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 7006 3340 7012 3392
rect 7064 3340 7070 3392
rect 7190 3340 7196 3392
rect 7248 3340 7254 3392
rect 1104 3290 11224 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 11224 3290
rect 1104 3216 11224 3238
rect 4154 3136 4160 3188
rect 4212 3136 4218 3188
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 5258 3176 5264 3188
rect 4387 3148 5264 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6086 3136 6092 3188
rect 6144 3176 6150 3188
rect 6457 3179 6515 3185
rect 6457 3176 6469 3179
rect 6144 3148 6469 3176
rect 6144 3136 6150 3148
rect 6457 3145 6469 3148
rect 6503 3145 6515 3179
rect 7098 3176 7104 3188
rect 6457 3139 6515 3145
rect 6840 3148 7104 3176
rect 3605 3111 3663 3117
rect 3605 3077 3617 3111
rect 3651 3108 3663 3111
rect 4172 3108 4200 3136
rect 4893 3111 4951 3117
rect 4893 3108 4905 3111
rect 3651 3080 3924 3108
rect 3651 3077 3663 3080
rect 3605 3071 3663 3077
rect 3510 3000 3516 3052
rect 3568 3000 3574 3052
rect 3786 3000 3792 3052
rect 3844 3000 3850 3052
rect 3896 3049 3924 3080
rect 4080 3080 4905 3108
rect 4080 3049 4108 3080
rect 4893 3077 4905 3080
rect 4939 3077 4951 3111
rect 4893 3071 4951 3077
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4246 3040 4252 3052
rect 4203 3012 4252 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3040 4583 3043
rect 4614 3040 4620 3052
rect 4571 3012 4620 3040
rect 4571 3009 4583 3012
rect 4525 3003 4583 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4798 3000 4804 3052
rect 4856 3000 4862 3052
rect 5166 3000 5172 3052
rect 5224 3000 5230 3052
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 5902 3040 5908 3052
rect 5307 3012 5908 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 5276 2972 5304 3003
rect 5902 3000 5908 3012
rect 5960 3000 5966 3052
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 6840 3040 6868 3148
rect 7098 3136 7104 3148
rect 7156 3176 7162 3188
rect 7156 3148 7604 3176
rect 7156 3136 7162 3148
rect 6914 3068 6920 3120
rect 6972 3108 6978 3120
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 6972 3080 7481 3108
rect 6972 3068 6978 3080
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 7576 3108 7604 3148
rect 7834 3136 7840 3188
rect 7892 3136 7898 3188
rect 8389 3111 8447 3117
rect 8389 3108 8401 3111
rect 7576 3080 8401 3108
rect 7469 3071 7527 3077
rect 8389 3077 8401 3080
rect 8435 3077 8447 3111
rect 8389 3071 8447 3077
rect 7008 3043 7066 3049
rect 7008 3040 7020 3043
rect 6840 3012 7020 3040
rect 7008 3009 7020 3012
rect 7054 3009 7066 3043
rect 7008 3003 7066 3009
rect 7101 3043 7159 3049
rect 7101 3009 7113 3043
rect 7147 3009 7159 3043
rect 7101 3003 7159 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 4764 2944 5304 2972
rect 4764 2932 4770 2944
rect 4522 2864 4528 2916
rect 4580 2904 4586 2916
rect 4617 2907 4675 2913
rect 4617 2904 4629 2907
rect 4580 2876 4629 2904
rect 4580 2864 4586 2876
rect 4617 2873 4629 2876
rect 4663 2873 4675 2907
rect 4617 2867 4675 2873
rect 6914 2796 6920 2848
rect 6972 2796 6978 2848
rect 7116 2836 7144 3003
rect 7208 2972 7236 3003
rect 7282 3000 7288 3052
rect 7340 3000 7346 3052
rect 7558 3000 7564 3052
rect 7616 3000 7622 3052
rect 7699 3043 7757 3049
rect 7699 3009 7711 3043
rect 7745 3040 7757 3043
rect 7926 3040 7932 3052
rect 7745 3012 7932 3040
rect 7745 3009 7757 3012
rect 7699 3003 7757 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 7374 2972 7380 2984
rect 7208 2944 7380 2972
rect 7374 2932 7380 2944
rect 7432 2972 7438 2984
rect 7432 2944 7972 2972
rect 7432 2932 7438 2944
rect 7944 2913 7972 2944
rect 7929 2907 7987 2913
rect 7929 2873 7941 2907
rect 7975 2873 7987 2907
rect 7929 2867 7987 2873
rect 8113 2907 8171 2913
rect 8113 2873 8125 2907
rect 8159 2873 8171 2907
rect 8113 2867 8171 2873
rect 8018 2836 8024 2848
rect 7116 2808 8024 2836
rect 8018 2796 8024 2808
rect 8076 2836 8082 2848
rect 8128 2836 8156 2867
rect 8076 2808 8156 2836
rect 8076 2796 8082 2808
rect 1104 2746 11224 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 11224 2746
rect 1104 2672 11224 2694
rect 3510 2592 3516 2644
rect 3568 2592 3574 2644
rect 4614 2592 4620 2644
rect 4672 2592 4678 2644
rect 5166 2592 5172 2644
rect 5224 2632 5230 2644
rect 5261 2635 5319 2641
rect 5261 2632 5273 2635
rect 5224 2604 5273 2632
rect 5224 2592 5230 2604
rect 5261 2601 5273 2604
rect 5307 2601 5319 2635
rect 5261 2595 5319 2601
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 6362 2632 6368 2644
rect 6227 2604 6368 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6362 2592 6368 2604
rect 6420 2592 6426 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7285 2635 7343 2641
rect 7285 2632 7297 2635
rect 7248 2604 7297 2632
rect 7248 2592 7254 2604
rect 7285 2601 7297 2604
rect 7331 2601 7343 2635
rect 7285 2595 7343 2601
rect 7558 2592 7564 2644
rect 7616 2632 7622 2644
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7616 2604 8033 2632
rect 7616 2592 7622 2604
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 8021 2595 8079 2601
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 8628 2604 8677 2632
rect 8628 2592 8634 2604
rect 8665 2601 8677 2604
rect 8711 2601 8723 2635
rect 8665 2595 8723 2601
rect 4157 2567 4215 2573
rect 4157 2533 4169 2567
rect 4203 2564 4215 2567
rect 4798 2564 4804 2576
rect 4203 2536 4804 2564
rect 4203 2533 4215 2536
rect 4157 2527 4215 2533
rect 4798 2524 4804 2536
rect 4856 2524 4862 2576
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 7377 2567 7435 2573
rect 7377 2564 7389 2567
rect 7064 2536 7389 2564
rect 7064 2524 7070 2536
rect 7377 2533 7389 2536
rect 7423 2533 7435 2567
rect 7377 2527 7435 2533
rect 6914 2456 6920 2508
rect 6972 2456 6978 2508
rect 7926 2496 7932 2508
rect 7668 2468 7932 2496
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 3329 2431 3387 2437
rect 3329 2428 3341 2431
rect 3292 2400 3341 2428
rect 3292 2388 3298 2400
rect 3329 2397 3341 2400
rect 3375 2397 3387 2431
rect 3329 2391 3387 2397
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3936 2400 3985 2428
rect 3936 2388 3942 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4580 2400 4813 2428
rect 4580 2388 4586 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5258 2388 5264 2440
rect 5316 2428 5322 2440
rect 5445 2431 5503 2437
rect 5445 2428 5457 2431
rect 5316 2400 5457 2428
rect 5316 2388 5322 2400
rect 5445 2397 5457 2400
rect 5491 2397 5503 2431
rect 5445 2391 5503 2397
rect 5997 2431 6055 2437
rect 5997 2397 6009 2431
rect 6043 2397 6055 2431
rect 5997 2391 6055 2397
rect 6012 2292 6040 2391
rect 6362 2388 6368 2440
rect 6420 2388 6426 2440
rect 6546 2437 6552 2440
rect 6519 2431 6552 2437
rect 6519 2397 6531 2431
rect 6519 2391 6552 2397
rect 6546 2388 6552 2391
rect 6604 2388 6610 2440
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6779 2400 7113 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 7101 2397 7113 2400
rect 7147 2428 7159 2431
rect 7282 2428 7288 2440
rect 7147 2400 7288 2428
rect 7147 2397 7159 2400
rect 7101 2391 7159 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7374 2388 7380 2440
rect 7432 2388 7438 2440
rect 7558 2388 7564 2440
rect 7616 2388 7622 2440
rect 7668 2437 7696 2468
rect 7926 2456 7932 2468
rect 7984 2456 7990 2508
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2397 7711 2431
rect 7653 2391 7711 2397
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 7760 2360 7788 2391
rect 7834 2388 7840 2440
rect 7892 2428 7898 2440
rect 8205 2431 8263 2437
rect 8205 2428 8217 2431
rect 7892 2400 8217 2428
rect 7892 2388 7898 2400
rect 8205 2397 8217 2400
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8481 2431 8539 2437
rect 8481 2428 8493 2431
rect 8444 2400 8493 2428
rect 8444 2388 8450 2400
rect 8481 2397 8493 2400
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 7484 2332 7788 2360
rect 6454 2292 6460 2304
rect 6012 2264 6460 2292
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7484 2292 7512 2332
rect 7156 2264 7512 2292
rect 7929 2295 7987 2301
rect 7156 2252 7162 2264
rect 7929 2261 7941 2295
rect 7975 2292 7987 2295
rect 8018 2292 8024 2304
rect 7975 2264 8024 2292
rect 7975 2261 7987 2264
rect 7929 2255 7987 2261
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 1104 2202 11224 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 11224 2202
rect 1104 2128 11224 2150
<< via1 >>
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 9404 11840 9456 11892
rect 4528 11772 4580 11824
rect 3884 11704 3936 11756
rect 4620 11568 4672 11620
rect 5264 11747 5316 11756
rect 5264 11713 5273 11747
rect 5273 11713 5307 11747
rect 5307 11713 5316 11747
rect 5264 11704 5316 11713
rect 5816 11704 5868 11756
rect 7104 11704 7156 11756
rect 7748 11704 7800 11756
rect 7932 11704 7984 11756
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 8484 11704 8536 11756
rect 9036 11704 9088 11756
rect 9128 11636 9180 11688
rect 6460 11568 6512 11620
rect 7564 11568 7616 11620
rect 8300 11568 8352 11620
rect 8944 11568 8996 11620
rect 5172 11500 5224 11552
rect 6276 11500 6328 11552
rect 7472 11500 7524 11552
rect 8484 11500 8536 11552
rect 9312 11500 9364 11552
rect 9496 11500 9548 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 7932 11339 7984 11348
rect 7932 11305 7941 11339
rect 7941 11305 7975 11339
rect 7975 11305 7984 11339
rect 7932 11296 7984 11305
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 5816 11228 5868 11280
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 5172 11135 5224 11144
rect 5172 11101 5181 11135
rect 5181 11101 5215 11135
rect 5215 11101 5224 11135
rect 5172 11092 5224 11101
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 6000 11092 6052 11144
rect 6276 11092 6328 11144
rect 6460 11135 6512 11144
rect 6460 11101 6469 11135
rect 6469 11101 6503 11135
rect 6503 11101 6512 11135
rect 6460 11092 6512 11101
rect 7380 11092 7432 11144
rect 8300 11160 8352 11212
rect 9128 11160 9180 11212
rect 4804 11067 4856 11076
rect 4804 11033 4813 11067
rect 4813 11033 4847 11067
rect 4847 11033 4856 11067
rect 4804 11024 4856 11033
rect 5632 11024 5684 11076
rect 7840 11024 7892 11076
rect 8116 11135 8168 11144
rect 8116 11101 8125 11135
rect 8125 11101 8159 11135
rect 8159 11101 8168 11135
rect 8116 11092 8168 11101
rect 8484 11135 8536 11144
rect 8484 11101 8492 11135
rect 8492 11101 8526 11135
rect 8526 11101 8536 11135
rect 8484 11092 8536 11101
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 9220 11092 9272 11144
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 9864 11135 9916 11144
rect 9864 11101 9877 11135
rect 9877 11101 9916 11135
rect 9496 11024 9548 11076
rect 9864 11092 9916 11101
rect 10876 11092 10928 11144
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 5908 10956 5960 11008
rect 7656 10956 7708 11008
rect 8300 10956 8352 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 3792 10752 3844 10804
rect 7656 10752 7708 10804
rect 4344 10684 4396 10736
rect 2964 10659 3016 10668
rect 2964 10625 2973 10659
rect 2973 10625 3007 10659
rect 3007 10625 3016 10659
rect 2964 10616 3016 10625
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 3792 10616 3844 10668
rect 4620 10616 4672 10668
rect 5632 10684 5684 10736
rect 7564 10684 7616 10736
rect 5172 10659 5224 10668
rect 5172 10625 5181 10659
rect 5181 10625 5215 10659
rect 5215 10625 5224 10659
rect 5172 10616 5224 10625
rect 5356 10616 5408 10668
rect 5724 10659 5776 10668
rect 5724 10625 5733 10659
rect 5733 10625 5767 10659
rect 5767 10625 5776 10659
rect 5724 10616 5776 10625
rect 7288 10616 7340 10668
rect 7748 10616 7800 10668
rect 2688 10548 2740 10600
rect 6828 10548 6880 10600
rect 6920 10591 6972 10600
rect 6920 10557 6929 10591
rect 6929 10557 6963 10591
rect 6963 10557 6972 10591
rect 6920 10548 6972 10557
rect 7840 10548 7892 10600
rect 8944 10659 8996 10668
rect 8944 10625 8953 10659
rect 8953 10625 8987 10659
rect 8987 10625 8996 10659
rect 8944 10616 8996 10625
rect 9220 10684 9272 10736
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 9588 10616 9640 10668
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 5080 10480 5132 10532
rect 7932 10480 7984 10532
rect 2136 10412 2188 10464
rect 3700 10455 3752 10464
rect 3700 10421 3709 10455
rect 3709 10421 3743 10455
rect 3743 10421 3752 10455
rect 3700 10412 3752 10421
rect 3884 10455 3936 10464
rect 3884 10421 3893 10455
rect 3893 10421 3927 10455
rect 3927 10421 3936 10455
rect 3884 10412 3936 10421
rect 6552 10412 6604 10464
rect 8760 10455 8812 10464
rect 8760 10421 8769 10455
rect 8769 10421 8803 10455
rect 8803 10421 8812 10455
rect 8760 10412 8812 10421
rect 9404 10412 9456 10464
rect 9772 10455 9824 10464
rect 9772 10421 9781 10455
rect 9781 10421 9815 10455
rect 9815 10421 9824 10455
rect 9772 10412 9824 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 3516 10208 3568 10260
rect 5080 10251 5132 10260
rect 5080 10217 5089 10251
rect 5089 10217 5123 10251
rect 5123 10217 5132 10251
rect 5080 10208 5132 10217
rect 6920 10208 6972 10260
rect 6552 10140 6604 10192
rect 7380 10208 7432 10260
rect 7932 10251 7984 10260
rect 7932 10217 7941 10251
rect 7941 10217 7975 10251
rect 7975 10217 7984 10251
rect 7932 10208 7984 10217
rect 7748 10140 7800 10192
rect 2136 10115 2188 10124
rect 2136 10081 2145 10115
rect 2145 10081 2179 10115
rect 2179 10081 2188 10115
rect 2136 10072 2188 10081
rect 4804 10072 4856 10124
rect 4160 10004 4212 10056
rect 5356 10004 5408 10056
rect 5816 10072 5868 10124
rect 6184 10115 6236 10124
rect 6184 10081 6193 10115
rect 6193 10081 6227 10115
rect 6227 10081 6236 10115
rect 6184 10072 6236 10081
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 2044 9936 2096 9988
rect 3884 9936 3936 9988
rect 6276 10047 6328 10056
rect 6276 10013 6285 10047
rect 6285 10013 6319 10047
rect 6319 10013 6328 10047
rect 6276 10004 6328 10013
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 6460 9936 6512 9988
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 8760 10208 8812 10260
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 9772 10072 9824 10124
rect 8208 10047 8260 10056
rect 8208 10013 8217 10047
rect 8217 10013 8251 10047
rect 8251 10013 8260 10047
rect 8208 10004 8260 10013
rect 9036 10004 9088 10056
rect 8300 9936 8352 9988
rect 10416 9936 10468 9988
rect 3976 9911 4028 9920
rect 3976 9877 3985 9911
rect 3985 9877 4019 9911
rect 4019 9877 4028 9911
rect 3976 9868 4028 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 8116 9664 8168 9716
rect 8208 9707 8260 9716
rect 8208 9673 8217 9707
rect 8217 9673 8251 9707
rect 8251 9673 8260 9707
rect 8208 9664 8260 9673
rect 9588 9664 9640 9716
rect 3700 9596 3752 9648
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 2780 9460 2832 9512
rect 4804 9528 4856 9580
rect 5540 9596 5592 9648
rect 5264 9528 5316 9580
rect 5816 9528 5868 9580
rect 8116 9571 8168 9580
rect 8116 9537 8125 9571
rect 8125 9537 8159 9571
rect 8159 9537 8168 9571
rect 8116 9528 8168 9537
rect 8576 9596 8628 9648
rect 10416 9596 10468 9648
rect 8392 9528 8444 9580
rect 9864 9528 9916 9580
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 4068 9460 4120 9512
rect 5724 9460 5776 9512
rect 9128 9460 9180 9512
rect 3884 9392 3936 9444
rect 4160 9392 4212 9444
rect 4620 9392 4672 9444
rect 5908 9392 5960 9444
rect 5632 9324 5684 9376
rect 6552 9324 6604 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 2780 9163 2832 9172
rect 2780 9129 2789 9163
rect 2789 9129 2823 9163
rect 2823 9129 2832 9163
rect 2780 9120 2832 9129
rect 4068 9120 4120 9172
rect 5448 9120 5500 9172
rect 5816 9163 5868 9172
rect 5816 9129 5825 9163
rect 5825 9129 5859 9163
rect 5859 9129 5868 9163
rect 5816 9120 5868 9129
rect 6368 9120 6420 9172
rect 3792 9052 3844 9104
rect 3976 8984 4028 9036
rect 4344 8916 4396 8968
rect 5264 9052 5316 9104
rect 5540 9052 5592 9104
rect 8208 9052 8260 9104
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 2964 8891 3016 8900
rect 2964 8857 2991 8891
rect 2991 8857 3016 8891
rect 2964 8848 3016 8857
rect 4068 8891 4120 8900
rect 4068 8857 4077 8891
rect 4077 8857 4111 8891
rect 4111 8857 4120 8891
rect 4068 8848 4120 8857
rect 8576 8984 8628 9036
rect 9036 9027 9088 9036
rect 9036 8993 9045 9027
rect 9045 8993 9079 9027
rect 9079 8993 9088 9027
rect 9036 8984 9088 8993
rect 9404 8984 9456 9036
rect 9956 8984 10008 9036
rect 4804 8848 4856 8900
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 6828 8916 6880 8968
rect 8116 8916 8168 8968
rect 8392 8959 8444 8968
rect 8392 8925 8401 8959
rect 8401 8925 8435 8959
rect 8435 8925 8444 8959
rect 8392 8916 8444 8925
rect 5540 8891 5592 8900
rect 5540 8857 5549 8891
rect 5549 8857 5583 8891
rect 5583 8857 5592 8891
rect 5540 8848 5592 8857
rect 6000 8891 6052 8900
rect 6000 8857 6009 8891
rect 6009 8857 6043 8891
rect 6043 8857 6052 8891
rect 6000 8848 6052 8857
rect 4436 8780 4488 8832
rect 4712 8780 4764 8832
rect 5816 8823 5868 8832
rect 5816 8789 5838 8823
rect 5838 8789 5868 8823
rect 5816 8780 5868 8789
rect 6184 8823 6236 8832
rect 6184 8789 6193 8823
rect 6193 8789 6227 8823
rect 6227 8789 6236 8823
rect 6184 8780 6236 8789
rect 6736 8848 6788 8900
rect 7196 8848 7248 8900
rect 9220 8848 9272 8900
rect 10324 8848 10376 8900
rect 6552 8780 6604 8832
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 9128 8780 9180 8832
rect 9680 8780 9732 8832
rect 9956 8780 10008 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5448 8576 5500 8628
rect 5540 8576 5592 8628
rect 6092 8576 6144 8628
rect 6644 8508 6696 8560
rect 3148 8440 3200 8492
rect 4528 8440 4580 8492
rect 1400 8372 1452 8424
rect 2044 8372 2096 8424
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 4620 8304 4672 8356
rect 5816 8440 5868 8492
rect 5448 8372 5500 8424
rect 5632 8372 5684 8424
rect 6276 8440 6328 8492
rect 8944 8576 8996 8628
rect 9128 8576 9180 8628
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 9312 8576 9364 8628
rect 7840 8508 7892 8560
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 10324 8619 10376 8628
rect 10324 8585 10333 8619
rect 10333 8585 10367 8619
rect 10367 8585 10376 8619
rect 10324 8576 10376 8585
rect 8852 8440 8904 8492
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 9404 8440 9456 8492
rect 9956 8440 10008 8492
rect 10232 8483 10284 8492
rect 10232 8449 10241 8483
rect 10241 8449 10275 8483
rect 10275 8449 10284 8483
rect 10232 8440 10284 8449
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 8116 8372 8168 8424
rect 6736 8304 6788 8356
rect 6828 8304 6880 8356
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 9634 8304 9686 8356
rect 10048 8304 10100 8356
rect 5724 8236 5776 8288
rect 6276 8236 6328 8288
rect 6368 8236 6420 8288
rect 7196 8236 7248 8288
rect 9220 8236 9272 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3148 8075 3200 8084
rect 3148 8041 3157 8075
rect 3157 8041 3191 8075
rect 3191 8041 3200 8075
rect 3148 8032 3200 8041
rect 6736 8075 6788 8084
rect 6736 8041 6745 8075
rect 6745 8041 6779 8075
rect 6779 8041 6788 8075
rect 6736 8032 6788 8041
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 7840 8032 7892 8084
rect 2688 7896 2740 7948
rect 3332 7896 3384 7948
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 6552 7964 6604 8016
rect 7104 7964 7156 8016
rect 3516 7896 3568 7948
rect 4160 7896 4212 7948
rect 5264 7939 5316 7948
rect 5264 7905 5273 7939
rect 5273 7905 5307 7939
rect 5307 7905 5316 7939
rect 5264 7896 5316 7905
rect 1584 7760 1636 7812
rect 3332 7760 3384 7812
rect 4712 7828 4764 7880
rect 4804 7828 4856 7880
rect 6368 7828 6420 7880
rect 8300 7896 8352 7948
rect 7840 7871 7892 7880
rect 7840 7837 7849 7871
rect 7849 7837 7883 7871
rect 7883 7837 7892 7871
rect 7840 7828 7892 7837
rect 5540 7760 5592 7812
rect 8024 7760 8076 7812
rect 3516 7692 3568 7744
rect 6184 7692 6236 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 3332 7531 3384 7540
rect 3332 7497 3341 7531
rect 3341 7497 3375 7531
rect 3375 7497 3384 7531
rect 3332 7488 3384 7497
rect 6000 7488 6052 7540
rect 9036 7488 9088 7540
rect 1492 7420 1544 7472
rect 3148 7395 3200 7404
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 4160 7420 4212 7472
rect 4620 7420 4672 7472
rect 6644 7420 6696 7472
rect 2688 7284 2740 7336
rect 1584 7216 1636 7268
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 9036 7352 9088 7404
rect 3516 7284 3568 7336
rect 3608 7216 3660 7268
rect 5816 7191 5868 7200
rect 5816 7157 5825 7191
rect 5825 7157 5859 7191
rect 5859 7157 5868 7191
rect 5816 7148 5868 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 6644 6987 6696 6996
rect 6644 6953 6653 6987
rect 6653 6953 6687 6987
rect 6687 6953 6696 6987
rect 6644 6944 6696 6953
rect 7196 6944 7248 6996
rect 1492 6808 1544 6860
rect 3700 6740 3752 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 7840 6740 7892 6792
rect 8944 6851 8996 6860
rect 8944 6817 8953 6851
rect 8953 6817 8987 6851
rect 8987 6817 8996 6851
rect 8944 6808 8996 6817
rect 10232 6808 10284 6860
rect 2044 6715 2096 6724
rect 2044 6681 2053 6715
rect 2053 6681 2087 6715
rect 2087 6681 2096 6715
rect 2044 6672 2096 6681
rect 9220 6715 9272 6724
rect 9220 6681 9229 6715
rect 9229 6681 9263 6715
rect 9263 6681 9272 6715
rect 9220 6672 9272 6681
rect 10232 6672 10284 6724
rect 2872 6604 2924 6656
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 7472 6604 7524 6656
rect 9496 6604 9548 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2044 6400 2096 6452
rect 7196 6400 7248 6452
rect 2872 6332 2924 6384
rect 3976 6332 4028 6384
rect 4620 6332 4672 6384
rect 6092 6375 6144 6384
rect 6092 6341 6101 6375
rect 6101 6341 6135 6375
rect 6135 6341 6144 6375
rect 6092 6332 6144 6341
rect 7472 6332 7524 6384
rect 8024 6400 8076 6452
rect 8852 6443 8904 6452
rect 8852 6409 8861 6443
rect 8861 6409 8895 6443
rect 8895 6409 8904 6443
rect 8852 6400 8904 6409
rect 9220 6400 9272 6452
rect 10232 6400 10284 6452
rect 1492 6264 1544 6316
rect 5172 6264 5224 6316
rect 6460 6264 6512 6316
rect 8944 6332 8996 6384
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8576 6307 8628 6316
rect 8576 6273 8585 6307
rect 8585 6273 8619 6307
rect 8619 6273 8628 6307
rect 8576 6264 8628 6273
rect 8668 6307 8720 6316
rect 8668 6273 8677 6307
rect 8677 6273 8711 6307
rect 8711 6273 8720 6307
rect 8668 6264 8720 6273
rect 8760 6264 8812 6316
rect 3056 6196 3108 6248
rect 3608 6196 3660 6248
rect 5356 6196 5408 6248
rect 6092 6196 6144 6248
rect 9496 6196 9548 6248
rect 10324 6264 10376 6316
rect 3608 6060 3660 6112
rect 3700 6060 3752 6112
rect 4712 6060 4764 6112
rect 5080 6060 5132 6112
rect 8852 6128 8904 6180
rect 6920 6060 6972 6112
rect 9312 6103 9364 6112
rect 9312 6069 9321 6103
rect 9321 6069 9355 6103
rect 9355 6069 9364 6103
rect 9312 6060 9364 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 3056 5899 3108 5908
rect 3056 5865 3065 5899
rect 3065 5865 3099 5899
rect 3099 5865 3108 5899
rect 3056 5856 3108 5865
rect 3976 5856 4028 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 5172 5856 5224 5908
rect 7380 5856 7432 5908
rect 7748 5856 7800 5908
rect 2872 5720 2924 5772
rect 2688 5652 2740 5704
rect 3700 5652 3752 5704
rect 3792 5652 3844 5704
rect 4252 5652 4304 5704
rect 4620 5720 4672 5772
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5080 5720 5132 5729
rect 5172 5720 5224 5772
rect 8024 5788 8076 5840
rect 8576 5856 8628 5908
rect 8484 5788 8536 5840
rect 8760 5856 8812 5908
rect 3424 5627 3476 5636
rect 3424 5593 3433 5627
rect 3433 5593 3467 5627
rect 3467 5593 3476 5627
rect 3424 5584 3476 5593
rect 6920 5652 6972 5704
rect 7104 5652 7156 5704
rect 5816 5584 5868 5636
rect 6460 5516 6512 5568
rect 8576 5652 8628 5704
rect 10324 5899 10376 5908
rect 10324 5865 10333 5899
rect 10333 5865 10367 5899
rect 10367 5865 10376 5899
rect 10324 5856 10376 5865
rect 8300 5584 8352 5636
rect 9312 5652 9364 5704
rect 10324 5652 10376 5704
rect 9036 5584 9088 5636
rect 10416 5584 10468 5636
rect 8760 5516 8812 5568
rect 9312 5559 9364 5568
rect 9312 5525 9321 5559
rect 9321 5525 9355 5559
rect 9355 5525 9364 5559
rect 9312 5516 9364 5525
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 4252 5355 4304 5364
rect 4252 5321 4261 5355
rect 4261 5321 4295 5355
rect 4295 5321 4304 5355
rect 4252 5312 4304 5321
rect 4712 5312 4764 5364
rect 8300 5312 8352 5364
rect 8668 5312 8720 5364
rect 3424 5244 3476 5296
rect 3792 5244 3844 5296
rect 5632 5244 5684 5296
rect 10416 5312 10468 5364
rect 2504 5108 2556 5160
rect 2688 5219 2740 5228
rect 2688 5185 2697 5219
rect 2697 5185 2731 5219
rect 2731 5185 2740 5219
rect 2688 5176 2740 5185
rect 2872 5219 2924 5228
rect 2872 5185 2881 5219
rect 2881 5185 2915 5219
rect 2915 5185 2924 5219
rect 2872 5176 2924 5185
rect 3976 5176 4028 5228
rect 8852 5287 8904 5296
rect 8852 5253 8861 5287
rect 8861 5253 8895 5287
rect 8895 5253 8904 5287
rect 8852 5244 8904 5253
rect 10048 5244 10100 5296
rect 7748 5219 7800 5228
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 8300 5176 8352 5228
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 8944 5176 8996 5228
rect 5540 5040 5592 5092
rect 1768 4972 1820 5024
rect 2320 5015 2372 5024
rect 2320 4981 2329 5015
rect 2329 4981 2363 5015
rect 2363 4981 2372 5015
rect 2320 4972 2372 4981
rect 8668 4972 8720 5024
rect 9128 4972 9180 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2504 4768 2556 4820
rect 8760 4768 8812 4820
rect 1492 4675 1544 4684
rect 1492 4641 1501 4675
rect 1501 4641 1535 4675
rect 1535 4641 1544 4675
rect 1492 4632 1544 4641
rect 4620 4632 4672 4684
rect 5632 4632 5684 4684
rect 3792 4564 3844 4616
rect 8944 4675 8996 4684
rect 8944 4641 8953 4675
rect 8953 4641 8987 4675
rect 8987 4641 8996 4675
rect 8944 4632 8996 4641
rect 9312 4632 9364 4684
rect 7748 4564 7800 4616
rect 1768 4539 1820 4548
rect 1768 4505 1777 4539
rect 1777 4505 1811 4539
rect 1811 4505 1820 4539
rect 1768 4496 1820 4505
rect 4712 4496 4764 4548
rect 5540 4428 5592 4480
rect 6000 4428 6052 4480
rect 8300 4428 8352 4480
rect 9956 4496 10008 4548
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 2320 4224 2372 4276
rect 2688 4224 2740 4276
rect 8852 4267 8904 4276
rect 8852 4233 8861 4267
rect 8861 4233 8895 4267
rect 8895 4233 8904 4267
rect 8852 4224 8904 4233
rect 10416 4224 10468 4276
rect 2504 4088 2556 4140
rect 4160 4088 4212 4140
rect 4804 4088 4856 4140
rect 5540 4156 5592 4208
rect 3792 4020 3844 4072
rect 3976 4020 4028 4072
rect 4712 3952 4764 4004
rect 4896 3952 4948 4004
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 5540 4020 5592 4072
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 7840 4088 7892 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8392 4088 8444 4140
rect 5724 3952 5776 4004
rect 7564 4020 7616 4072
rect 8576 4020 8628 4072
rect 9128 4131 9180 4140
rect 9128 4097 9137 4131
rect 9137 4097 9171 4131
rect 9171 4097 9180 4131
rect 9128 4088 9180 4097
rect 9956 4088 10008 4140
rect 10324 4088 10376 4140
rect 10876 4131 10928 4140
rect 10876 4097 10885 4131
rect 10885 4097 10919 4131
rect 10919 4097 10928 4131
rect 10876 4088 10928 4097
rect 5356 3884 5408 3936
rect 7288 3884 7340 3936
rect 7932 3884 7984 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 2504 3680 2556 3732
rect 4160 3680 4212 3732
rect 4804 3680 4856 3732
rect 5540 3723 5592 3732
rect 5540 3689 5549 3723
rect 5549 3689 5583 3723
rect 5583 3689 5592 3723
rect 5540 3680 5592 3689
rect 6552 3680 6604 3732
rect 7380 3680 7432 3732
rect 8576 3680 8628 3732
rect 4068 3519 4120 3528
rect 4068 3485 4077 3519
rect 4077 3485 4111 3519
rect 4111 3485 4120 3519
rect 4068 3476 4120 3485
rect 4160 3519 4212 3528
rect 4160 3485 4169 3519
rect 4169 3485 4203 3519
rect 4203 3485 4212 3519
rect 4160 3476 4212 3485
rect 4896 3476 4948 3528
rect 6000 3587 6052 3596
rect 6000 3553 6009 3587
rect 6009 3553 6043 3587
rect 6043 3553 6052 3587
rect 6000 3544 6052 3553
rect 4528 3408 4580 3460
rect 4712 3451 4764 3460
rect 4712 3417 4721 3451
rect 4721 3417 4755 3451
rect 4755 3417 4764 3451
rect 4712 3408 4764 3417
rect 5724 3519 5776 3528
rect 5724 3485 5733 3519
rect 5733 3485 5767 3519
rect 5767 3485 5776 3519
rect 5724 3476 5776 3485
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 6092 3519 6144 3528
rect 6092 3485 6101 3519
rect 6101 3485 6135 3519
rect 6135 3485 6144 3519
rect 6092 3476 6144 3485
rect 6552 3476 6604 3528
rect 7564 3612 7616 3664
rect 7564 3476 7616 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8576 3519 8628 3528
rect 8576 3485 8584 3519
rect 8584 3485 8618 3519
rect 8618 3485 8628 3519
rect 8576 3476 8628 3485
rect 9128 3476 9180 3528
rect 5264 3340 5316 3392
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 4160 3136 4212 3188
rect 5264 3136 5316 3188
rect 6092 3136 6144 3188
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 4252 3000 4304 3052
rect 4620 3000 4672 3052
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 4804 3000 4856 3009
rect 5172 3043 5224 3052
rect 5172 3009 5181 3043
rect 5181 3009 5215 3043
rect 5215 3009 5224 3043
rect 5172 3000 5224 3009
rect 4712 2932 4764 2984
rect 5908 3000 5960 3052
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7104 3136 7156 3188
rect 6920 3068 6972 3120
rect 7840 3179 7892 3188
rect 7840 3145 7849 3179
rect 7849 3145 7883 3179
rect 7883 3145 7892 3179
rect 7840 3136 7892 3145
rect 4528 2864 4580 2916
rect 6920 2839 6972 2848
rect 6920 2805 6929 2839
rect 6929 2805 6963 2839
rect 6963 2805 6972 2839
rect 6920 2796 6972 2805
rect 7288 3043 7340 3052
rect 7288 3009 7298 3043
rect 7298 3009 7332 3043
rect 7332 3009 7340 3043
rect 7288 3000 7340 3009
rect 7564 3043 7616 3052
rect 7564 3009 7573 3043
rect 7573 3009 7607 3043
rect 7607 3009 7616 3043
rect 7564 3000 7616 3009
rect 7932 3000 7984 3052
rect 7380 2932 7432 2984
rect 8024 2796 8076 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 3516 2635 3568 2644
rect 3516 2601 3525 2635
rect 3525 2601 3559 2635
rect 3559 2601 3568 2635
rect 3516 2592 3568 2601
rect 4620 2635 4672 2644
rect 4620 2601 4629 2635
rect 4629 2601 4663 2635
rect 4663 2601 4672 2635
rect 4620 2592 4672 2601
rect 5172 2592 5224 2644
rect 6368 2592 6420 2644
rect 7196 2592 7248 2644
rect 7564 2592 7616 2644
rect 8576 2592 8628 2644
rect 4804 2524 4856 2576
rect 7012 2524 7064 2576
rect 6920 2499 6972 2508
rect 6920 2465 6929 2499
rect 6929 2465 6963 2499
rect 6963 2465 6972 2499
rect 6920 2456 6972 2465
rect 3240 2388 3292 2440
rect 3884 2388 3936 2440
rect 4528 2388 4580 2440
rect 5264 2388 5316 2440
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 6552 2431 6604 2440
rect 6552 2397 6565 2431
rect 6565 2397 6604 2431
rect 6552 2388 6604 2397
rect 7288 2388 7340 2440
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 7564 2431 7616 2440
rect 7564 2397 7573 2431
rect 7573 2397 7607 2431
rect 7607 2397 7616 2431
rect 7564 2388 7616 2397
rect 7932 2456 7984 2508
rect 7840 2388 7892 2440
rect 8392 2388 8444 2440
rect 6460 2252 6512 2304
rect 7104 2252 7156 2304
rect 8024 2252 8076 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 3882 13716 3938 14516
rect 4526 13716 4582 14516
rect 5170 13716 5226 14516
rect 5814 13716 5870 14516
rect 7102 13716 7158 14516
rect 7746 13716 7802 14516
rect 8390 13716 8446 14516
rect 9034 13716 9090 14516
rect 3896 11762 3924 13716
rect 4540 11830 4568 13716
rect 5184 12730 5212 13716
rect 5184 12702 5304 12730
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 5276 11762 5304 12702
rect 5828 11762 5856 13716
rect 7116 11762 7144 13716
rect 7760 11762 7788 13716
rect 8404 12434 8432 13716
rect 8404 12406 8524 12434
rect 8496 11762 8524 12406
rect 9048 11762 9076 13716
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 7748 11756 7800 11762
rect 7748 11698 7800 11704
rect 7932 11756 7984 11762
rect 7932 11698 7984 11704
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10810 3832 10950
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 4356 10742 4384 11086
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4632 10674 4660 11562
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 6276 11552 6328 11558
rect 6276 11494 6328 11500
rect 5184 11150 5212 11494
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5172 11144 5224 11150
rect 5356 11144 5408 11150
rect 5224 11092 5304 11098
rect 5172 11086 5304 11092
rect 5356 11086 5408 11092
rect 4804 11076 4856 11082
rect 5184 11070 5304 11086
rect 4804 11018 4856 11024
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3792 10668 3844 10674
rect 3792 10610 3844 10616
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2136 10464 2188 10470
rect 2136 10406 2188 10412
rect 2148 10130 2176 10406
rect 2136 10124 2188 10130
rect 2136 10066 2188 10072
rect 2044 9988 2096 9994
rect 2044 9930 2096 9936
rect 2056 9518 2084 9930
rect 2044 9512 2096 9518
rect 2044 9454 2096 9460
rect 2056 8430 2084 9454
rect 1400 8424 1452 8430
rect 1400 8366 1452 8372
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 1412 7886 1440 8366
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7426 1440 7822
rect 1504 7585 1532 8298
rect 2700 7954 2728 10542
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 9178 2820 9454
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2976 8906 3004 10610
rect 3528 10266 3556 10610
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3712 9654 3740 10406
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3804 9110 3832 10610
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 9994 3924 10406
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3884 9988 3936 9994
rect 3884 9930 3936 9936
rect 3976 9920 4028 9926
rect 3976 9862 4028 9868
rect 3884 9444 3936 9450
rect 3884 9386 3936 9392
rect 3792 9104 3844 9110
rect 3792 9046 3844 9052
rect 2964 8900 3016 8906
rect 2964 8842 3016 8848
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3160 8090 3188 8434
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 2688 7948 2740 7954
rect 2688 7890 2740 7896
rect 1584 7812 1636 7818
rect 1584 7754 1636 7760
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 1492 7472 1544 7478
rect 1412 7420 1492 7426
rect 1412 7414 1544 7420
rect 1412 7398 1532 7414
rect 1504 6866 1532 7398
rect 1596 7274 1624 7754
rect 2700 7342 2728 7890
rect 3160 7410 3188 8026
rect 3332 7948 3384 7954
rect 3516 7948 3568 7954
rect 3384 7908 3516 7936
rect 3332 7890 3384 7896
rect 3332 7812 3384 7818
rect 3332 7754 3384 7760
rect 3344 7546 3372 7754
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 3148 7404 3200 7410
rect 3148 7346 3200 7352
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 1584 7268 1636 7274
rect 1584 7210 1636 7216
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 6322 1532 6802
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2056 6458 2084 6666
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2884 6390 2912 6598
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1504 4690 1532 6258
rect 2884 5778 2912 6326
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3068 5914 3096 6190
rect 3056 5908 3108 5914
rect 3056 5850 3108 5856
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2700 5234 2728 5646
rect 2884 5234 2912 5714
rect 3436 5642 3464 7908
rect 3516 7890 3568 7896
rect 3516 7744 3568 7750
rect 3516 7686 3568 7692
rect 3528 7342 3556 7686
rect 3804 7426 3832 9046
rect 3896 8922 3924 9386
rect 3988 9042 4016 9862
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 9178 4108 9454
rect 4172 9450 4200 9998
rect 4632 9450 4660 10610
rect 4816 10130 4844 11018
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 5276 10690 5304 11070
rect 5184 10674 5304 10690
rect 5368 10674 5396 11086
rect 5632 11076 5684 11082
rect 5632 11018 5684 11024
rect 5644 10742 5672 11018
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5172 10668 5304 10674
rect 5224 10662 5304 10668
rect 5356 10668 5408 10674
rect 5172 10610 5224 10616
rect 5356 10610 5408 10616
rect 5080 10532 5132 10538
rect 5080 10474 5132 10480
rect 5092 10266 5120 10474
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4804 10124 4856 10130
rect 4804 10066 4856 10072
rect 4816 9586 4844 10066
rect 5092 10010 5120 10202
rect 5368 10062 5396 10610
rect 5356 10056 5408 10062
rect 5092 9982 5304 10010
rect 5356 9998 5408 10004
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5276 9586 5304 9982
rect 5552 9654 5580 9998
rect 5540 9648 5592 9654
rect 5354 9616 5410 9625
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 5264 9580 5316 9586
rect 5540 9590 5592 9596
rect 5354 9551 5410 9560
rect 5264 9522 5316 9528
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4620 9444 4672 9450
rect 4620 9386 4672 9392
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 5264 9104 5316 9110
rect 5264 9046 5316 9052
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4344 8968 4396 8974
rect 3896 8906 4108 8922
rect 4528 8968 4580 8974
rect 4396 8916 4476 8922
rect 4344 8910 4476 8916
rect 4528 8910 4580 8916
rect 3896 8900 4120 8906
rect 3896 8894 4068 8900
rect 4356 8894 4476 8910
rect 4068 8842 4120 8848
rect 4448 8838 4476 8894
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4540 8498 4568 8910
rect 4804 8900 4856 8906
rect 4804 8842 4856 8848
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4160 7948 4212 7954
rect 4160 7890 4212 7896
rect 4172 7478 4200 7890
rect 4632 7478 4660 8298
rect 4724 7886 4752 8774
rect 4816 7886 4844 8842
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 7954 5304 9046
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 3712 7398 3832 7426
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4620 7472 4672 7478
rect 4620 7414 4672 7420
rect 3516 7336 3568 7342
rect 3712 7290 3740 7398
rect 3516 7278 3568 7284
rect 3620 7274 3740 7290
rect 3608 7268 3740 7274
rect 3660 7262 3740 7268
rect 3608 7210 3660 7216
rect 3712 6798 3740 7262
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 5368 6798 5396 9551
rect 5644 9382 5672 10678
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5736 9518 5764 10610
rect 5828 10130 5856 11222
rect 6288 11150 6316 11494
rect 6472 11150 6500 11562
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11234 7512 11494
rect 7392 11206 7512 11234
rect 7392 11150 7420 11206
rect 6000 11144 6052 11150
rect 6276 11144 6328 11150
rect 6052 11092 6224 11098
rect 6000 11086 6224 11092
rect 6276 11086 6328 11092
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 6012 11070 6224 11086
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5920 10062 5948 10950
rect 6196 10130 6224 11070
rect 6184 10124 6236 10130
rect 6184 10066 6236 10072
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5632 9376 5684 9382
rect 5632 9318 5684 9324
rect 5828 9178 5856 9522
rect 5920 9450 5948 9998
rect 5908 9444 5960 9450
rect 5908 9386 5960 9392
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5816 9172 5868 9178
rect 5816 9114 5868 9120
rect 5460 8634 5488 9114
rect 5540 9104 5592 9110
rect 5540 9046 5592 9052
rect 5552 8906 5580 9046
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5552 8634 5580 8842
rect 5816 8832 5868 8838
rect 5816 8774 5868 8780
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5552 8514 5580 8570
rect 5460 8486 5580 8514
rect 5828 8498 5856 8774
rect 5816 8492 5868 8498
rect 5460 8430 5488 8486
rect 5816 8434 5868 8440
rect 5448 8424 5500 8430
rect 5632 8424 5684 8430
rect 5448 8366 5500 8372
rect 5552 8372 5632 8378
rect 5552 8366 5684 8372
rect 5552 8350 5672 8366
rect 5552 7818 5580 8350
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5736 7410 5764 8230
rect 6012 7546 6040 8842
rect 6196 8838 6224 10066
rect 6288 10062 6316 11086
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6472 9994 6500 11086
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6920 10600 6972 10606
rect 6920 10542 6972 10548
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 10198 6592 10406
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6564 10062 6592 10134
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6460 9988 6512 9994
rect 6460 9930 6512 9936
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6380 8974 6408 9114
rect 6564 8974 6592 9318
rect 6840 8974 6868 10542
rect 6932 10266 6960 10542
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6564 8838 6592 8910
rect 6736 8900 6788 8906
rect 6736 8842 6788 8848
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6092 8628 6144 8634
rect 6092 8570 6144 8576
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3712 6202 3740 6734
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 4620 6384 4672 6390
rect 4620 6326 4672 6332
rect 3620 6118 3648 6190
rect 3712 6174 3832 6202
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3700 6112 3752 6118
rect 3700 6054 3752 6060
rect 3712 5710 3740 6054
rect 3804 5710 3832 6174
rect 3988 5914 4016 6326
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5914 4660 6326
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3436 5302 3464 5578
rect 3804 5302 3832 5646
rect 4264 5370 4292 5646
rect 4252 5364 4304 5370
rect 4252 5306 4304 5312
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 1492 4684 1544 4690
rect 1492 4626 1544 4632
rect 1780 4554 1808 4966
rect 1768 4548 1820 4554
rect 1768 4490 1820 4496
rect 2332 4282 2360 4966
rect 2516 4826 2544 5102
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2516 4146 2544 4762
rect 2700 4282 2728 5170
rect 3804 4622 3832 5238
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2516 3738 2544 4082
rect 3988 4078 4016 5170
rect 4264 5012 4292 5306
rect 4080 4984 4292 5012
rect 4080 4808 4108 4984
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4080 4780 4200 4808
rect 4172 4146 4200 4780
rect 4632 4690 4660 5714
rect 4724 5370 4752 6054
rect 5092 5778 5120 6054
rect 5184 5914 5212 6258
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5184 5778 5212 5850
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 5172 5772 5224 5778
rect 5172 5714 5224 5720
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4724 4706 4752 5306
rect 4620 4684 4672 4690
rect 4724 4678 4844 4706
rect 4620 4626 4672 4632
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 3804 3058 3832 4014
rect 4724 4010 4752 4490
rect 4816 4146 4844 4678
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4712 4004 4764 4010
rect 4712 3946 4764 3952
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4816 3738 4844 4082
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4172 3618 4200 3674
rect 4080 3590 4292 3618
rect 4080 3534 4108 3590
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4172 3194 4200 3470
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4264 3058 4292 3590
rect 4908 3534 4936 3946
rect 5368 3942 5396 6190
rect 5828 5642 5856 7142
rect 6104 6390 6132 8570
rect 6196 7750 6224 8774
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6288 8294 6316 8434
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6380 7886 6408 8230
rect 6564 8022 6592 8774
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6184 7744 6236 7750
rect 6184 7686 6236 7692
rect 6656 7478 6684 8502
rect 6748 8362 6776 8842
rect 6840 8362 6868 8910
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6748 8090 6776 8298
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 7116 8022 7144 8366
rect 7208 8294 7236 8842
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 8090 7236 8230
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6656 7002 6684 7414
rect 7208 7002 7236 8026
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7208 6458 7236 6598
rect 7196 6452 7248 6458
rect 7196 6394 7248 6400
rect 6092 6384 6144 6390
rect 6092 6326 6144 6332
rect 6104 6254 6132 6326
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 6472 5574 6500 6258
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5710 6960 6054
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5552 4486 5580 5034
rect 5644 4690 5672 5238
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5552 4214 5580 4422
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5552 3738 5580 4014
rect 5724 4004 5776 4010
rect 5724 3946 5776 3952
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5736 3534 5764 3946
rect 6012 3602 6040 4422
rect 6472 3618 6500 5510
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6564 3738 6592 4082
rect 6552 3732 6604 3738
rect 6552 3674 6604 3680
rect 6000 3596 6052 3602
rect 6472 3590 6592 3618
rect 6000 3538 6052 3544
rect 6564 3534 6592 3590
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 4528 3460 4580 3466
rect 4528 3402 4580 3408
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 3528 2650 3556 2994
rect 4540 2922 4568 3402
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4528 2916 4580 2922
rect 4528 2858 4580 2864
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 2994
rect 4724 2990 4752 3402
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 5276 3194 5304 3334
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5920 3058 5948 3470
rect 6104 3194 6132 3470
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6368 3052 6420 3058
rect 6368 2994 6420 3000
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4816 2582 4844 2994
rect 5184 2650 5212 2994
rect 6380 2650 6408 2994
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 6368 2644 6420 2650
rect 6368 2586 6420 2592
rect 4804 2576 4856 2582
rect 4804 2518 4856 2524
rect 6380 2446 6408 2586
rect 6564 2446 6592 3470
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 6932 2854 6960 3062
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2514 6960 2790
rect 7024 2582 7052 3334
rect 7116 3194 7144 5646
rect 7300 3942 7328 10610
rect 7392 10266 7420 11086
rect 7576 10742 7604 11562
rect 7944 11354 7972 11698
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 8312 11218 8340 11562
rect 8404 11354 8432 11698
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 8944 11620 8996 11626
rect 8944 11562 8996 11568
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8496 11150 8524 11494
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 10810 7696 10950
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7576 10062 7604 10678
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7668 8090 7696 10746
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7760 10198 7788 10610
rect 7852 10606 7880 11018
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7932 10532 7984 10538
rect 7932 10474 7984 10480
rect 7944 10266 7972 10474
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7748 10192 7800 10198
rect 7748 10134 7800 10140
rect 8128 9722 8156 11086
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8220 9722 8248 9998
rect 8312 9994 8340 10950
rect 8300 9988 8352 9994
rect 8300 9930 8352 9936
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8128 8974 8156 9522
rect 8220 9110 8248 9658
rect 8588 9654 8616 11086
rect 8956 10674 8984 11562
rect 9140 11218 9168 11630
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9232 10742 9260 11086
rect 9220 10736 9272 10742
rect 9220 10678 9272 10684
rect 9324 10674 9352 11494
rect 9416 11150 9444 11834
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9416 10470 9444 11086
rect 9508 11082 9536 11494
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 8772 10266 8800 10406
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 9036 10056 9088 10062
rect 9036 9998 9088 10004
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8208 9104 8260 9110
rect 8208 9046 8260 9052
rect 8404 8974 8432 9522
rect 8588 9042 8616 9590
rect 9048 9042 9076 9998
rect 9600 9722 9628 10610
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10130 9812 10406
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 9876 9586 9904 11086
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 8116 8968 8168 8974
rect 8116 8910 8168 8916
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7852 8090 7880 8502
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7840 8084 7892 8090
rect 7840 8026 7892 8032
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 6798 7880 7822
rect 8036 7818 8064 8774
rect 8128 8430 8156 8910
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 8588 8362 8616 8978
rect 9048 8650 9076 8978
rect 9140 8838 9168 9454
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9956 9036 10008 9042
rect 9956 8978 10008 8984
rect 9220 8900 9272 8906
rect 9220 8842 9272 8848
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8956 8634 9076 8650
rect 9140 8634 9168 8774
rect 9232 8634 9260 8842
rect 8944 8628 9076 8634
rect 8996 8622 9076 8628
rect 8944 8570 8996 8576
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7392 5914 7420 6598
rect 7484 6390 7512 6598
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7760 5914 7788 6734
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 7760 5234 7788 5850
rect 8036 5846 8064 6394
rect 8312 6322 8340 7890
rect 8864 6458 8892 8434
rect 9048 7546 9076 8622
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9324 8498 9352 8570
rect 9416 8498 9444 8978
rect 9968 8838 9996 8978
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 9692 8634 9720 8774
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9968 8498 9996 8774
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 9218 8392 9274 8401
rect 9218 8327 9274 8336
rect 9586 8392 9642 8401
rect 9642 8362 9674 8378
rect 10060 8362 10088 10610
rect 10888 10266 10916 11086
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10416 9988 10468 9994
rect 10416 9930 10468 9936
rect 10428 9654 10456 9930
rect 10416 9648 10468 9654
rect 10416 9590 10468 9596
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 8498 10272 9522
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 8634 10364 8842
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 9642 8356 9686 8362
rect 9586 8327 9634 8336
rect 9232 8294 9260 8327
rect 9634 8298 9686 8304
rect 10048 8356 10100 8362
rect 10048 8298 10100 8304
rect 9220 8288 9272 8294
rect 9272 8248 9352 8276
rect 9220 8230 9272 8236
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9048 7410 9076 7482
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9048 7154 9076 7346
rect 8956 7126 9076 7154
rect 8956 6866 8984 7126
rect 8944 6860 8996 6866
rect 8944 6802 8996 6808
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8668 6316 8720 6322
rect 8668 6258 8720 6264
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8588 5914 8616 6258
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8024 5840 8076 5846
rect 8024 5782 8076 5788
rect 8484 5840 8536 5846
rect 8484 5782 8536 5788
rect 8300 5636 8352 5642
rect 8300 5578 8352 5584
rect 8312 5386 8340 5578
rect 8312 5370 8432 5386
rect 8300 5364 8432 5370
rect 8352 5358 8432 5364
rect 8300 5306 8352 5312
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7760 4622 7788 5170
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 8312 4486 8340 5170
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4146 8340 4422
rect 8404 4146 8432 5358
rect 8496 5234 8524 5782
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7392 3738 7420 4082
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7576 3670 7604 4014
rect 7564 3664 7616 3670
rect 7564 3606 7616 3612
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 7208 2650 7236 3334
rect 7576 3058 7604 3470
rect 7852 3194 7880 4082
rect 8588 4078 8616 5646
rect 8680 5370 8708 6258
rect 8772 5914 8800 6258
rect 8864 6186 8892 6394
rect 8956 6390 8984 6802
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9232 6458 9260 6666
rect 9220 6452 9272 6458
rect 9220 6394 9272 6400
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8666 5128 8722 5137
rect 8666 5063 8722 5072
rect 8680 5030 8708 5063
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8772 4826 8800 5510
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8864 4282 8892 5238
rect 8956 5234 8984 6326
rect 9324 6118 9352 8248
rect 10244 6882 10272 8434
rect 10244 6866 10364 6882
rect 10232 6860 10364 6866
rect 10284 6854 10364 6860
rect 10232 6802 10284 6808
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9508 6254 9536 6598
rect 10244 6458 10272 6666
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10336 6322 10364 6854
rect 10324 6316 10376 6322
rect 10324 6258 10376 6264
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9324 5710 9352 6054
rect 10336 5914 10364 6258
rect 10324 5908 10376 5914
rect 10324 5850 10376 5856
rect 10336 5710 10364 5850
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 4690 8984 5170
rect 9048 5137 9076 5578
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9034 5128 9090 5137
rect 9034 5063 9090 5072
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 9140 4146 9168 4966
rect 9324 4690 9352 5510
rect 10060 5302 10088 5510
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9968 4146 9996 4490
rect 10336 4146 10364 5646
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10428 5370 10456 5578
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10428 4282 10456 5306
rect 10874 4856 10930 4865
rect 10874 4791 10930 4800
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10888 4146 10916 4791
rect 9128 4140 9180 4146
rect 9128 4082 9180 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7944 3534 7972 3878
rect 8588 3738 8616 4014
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 9140 3534 9168 4082
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7944 3058 7972 3470
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7300 2446 7328 2994
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7392 2446 7420 2926
rect 7576 2650 7604 2994
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7576 2446 7604 2586
rect 7944 2514 7972 2994
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7564 2440 7616 2446
rect 7840 2440 7892 2446
rect 7564 2382 7616 2388
rect 7760 2400 7840 2428
rect 3252 800 3280 2382
rect 3896 800 3924 2382
rect 4540 800 4568 2382
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1306 5304 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 5184 1278 5304 1306
rect 5184 800 5212 1278
rect 6472 800 6500 2246
rect 7116 800 7144 2246
rect 7760 800 7788 2400
rect 7840 2382 7892 2388
rect 8036 2310 8064 2790
rect 8588 2650 8616 3470
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8404 800 8432 2382
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
<< via2 >>
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 1490 7520 1546 7576
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5354 9560 5410 9616
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 9218 8336 9274 8392
rect 9586 8356 9642 8392
rect 9586 8336 9634 8356
rect 9634 8336 9642 8356
rect 8666 5072 8722 5128
rect 9034 5072 9090 5128
rect 10874 4800 10930 4856
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
<< metal3 >>
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 5349 9618 5415 9621
rect 0 9616 5415 9618
rect 0 9560 5354 9616
rect 5410 9560 5415 9616
rect 0 9558 5415 9560
rect 0 9528 800 9558
rect 5349 9555 5415 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 9213 8394 9279 8397
rect 9581 8394 9647 8397
rect 9213 8392 9647 8394
rect 9213 8336 9218 8392
rect 9274 8336 9586 8392
rect 9642 8336 9647 8392
rect 9213 8334 9647 8336
rect 9213 8331 9279 8334
rect 9581 8331 9647 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1485 7578 1551 7581
rect 0 7576 1551 7578
rect 0 7520 1490 7576
rect 1546 7520 1551 7576
rect 0 7518 1551 7520
rect 0 7488 800 7518
rect 1485 7515 1551 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 8661 5130 8727 5133
rect 9029 5130 9095 5133
rect 8661 5128 9095 5130
rect 8661 5072 8666 5128
rect 8722 5072 9034 5128
rect 9090 5072 9095 5128
rect 8661 5070 9095 5072
rect 8661 5067 8727 5070
rect 9029 5067 9095 5070
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 10869 4858 10935 4861
rect 11572 4858 12372 4888
rect 10869 4856 12372 4858
rect 10869 4800 10874 4856
rect 10930 4800 12372 4856
rect 10869 4798 12372 4800
rect 10869 4795 10935 4798
rect 11572 4768 12372 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 11456 4528 12016
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 12000 5188 12016
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _113_
timestamp 0
transform -1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _114_
timestamp 0
transform -1 0 4692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _115_
timestamp 0
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_
timestamp 0
transform 1 0 5428 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _117_
timestamp 0
transform -1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 0
transform -1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 0
transform -1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 0
transform -1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _121_
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 0
transform 1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _123_
timestamp 0
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 0
transform 1 0 4784 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _125_
timestamp 0
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126_
timestamp 0
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _127_
timestamp 0
transform -1 0 5520 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _128_
timestamp 0
transform -1 0 6164 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _129_
timestamp 0
transform 1 0 4048 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _130_
timestamp 0
transform 1 0 5704 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _131_
timestamp 0
transform -1 0 5428 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _132_
timestamp 0
transform 1 0 5704 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _133_
timestamp 0
transform 1 0 6164 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or4bb_4  _134_
timestamp 0
transform -1 0 5704 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2b_1  _135_
timestamp 0
transform 1 0 9660 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _136_
timestamp 0
transform 1 0 9292 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _137_
timestamp 0
transform -1 0 8648 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _138_
timestamp 0
transform 1 0 7544 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _139_
timestamp 0
transform -1 0 8188 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand4_1  _140_
timestamp 0
transform 1 0 8280 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _141_
timestamp 0
transform -1 0 9292 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _142_
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _143_
timestamp 0
transform 1 0 6900 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _144_
timestamp 0
transform 1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _145_
timestamp 0
transform -1 0 4416 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _146_
timestamp 0
transform -1 0 4416 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _147_
timestamp 0
transform -1 0 5612 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _148_
timestamp 0
transform -1 0 8740 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _149_
timestamp 0
transform 1 0 5704 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _150_
timestamp 0
transform -1 0 7176 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _151_
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _152_
timestamp 0
transform 1 0 6900 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _153_
timestamp 0
transform 1 0 7636 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _154_
timestamp 0
transform -1 0 8464 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _155_
timestamp 0
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _156_
timestamp 0
transform -1 0 7452 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _157_
timestamp 0
transform 1 0 7176 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _158_
timestamp 0
transform 1 0 6992 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _159_
timestamp 0
transform -1 0 6900 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _160_
timestamp 0
transform 1 0 6992 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _161_
timestamp 0
transform -1 0 6808 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_4  _162_
timestamp 0
transform -1 0 8648 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__o211a_4  _163_
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1326 592
use sky130_fd_sc_hd__xnor2_1  _164_
timestamp 0
transform -1 0 2024 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _165_
timestamp 0
transform -1 0 2668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _166_
timestamp 0
transform 1 0 2576 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _167_
timestamp 0
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _168_
timestamp 0
transform -1 0 3496 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _169_
timestamp 0
transform 1 0 2392 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _170_
timestamp 0
transform -1 0 2944 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 0
transform -1 0 2576 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _172_
timestamp 0
transform 1 0 4876 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _173_
timestamp 0
transform -1 0 4876 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _174_
timestamp 0
transform 1 0 4232 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _175_
timestamp 0
transform 1 0 5244 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _176_
timestamp 0
transform 1 0 4508 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _177_
timestamp 0
transform -1 0 6164 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _178_
timestamp 0
transform -1 0 7268 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _179_
timestamp 0
transform 1 0 7728 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _180_
timestamp 0
transform 1 0 7268 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _181_
timestamp 0
transform -1 0 7820 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _182_
timestamp 0
transform 1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _183_
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _184_
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _185_
timestamp 0
transform 1 0 8648 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _186_
timestamp 0
transform 1 0 8004 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _187_
timestamp 0
transform -1 0 8740 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _188_
timestamp 0
transform 1 0 8464 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _189_
timestamp 0
transform 1 0 9568 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _190_
timestamp 0
transform 1 0 8280 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _191_
timestamp 0
transform 1 0 8924 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _192_
timestamp 0
transform 1 0 9568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _193_
timestamp 0
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _194_
timestamp 0
transform 1 0 8648 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _195_
timestamp 0
transform 1 0 8648 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _196_
timestamp 0
transform -1 0 10212 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _197_
timestamp 0
transform 1 0 8004 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _198_
timestamp 0
transform -1 0 8556 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _199_
timestamp 0
transform 1 0 6808 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _200_
timestamp 0
transform -1 0 5428 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _201_
timestamp 0
transform -1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _202_
timestamp 0
transform -1 0 5612 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _203_
timestamp 0
transform -1 0 6072 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _204_
timestamp 0
transform 1 0 4600 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _205_
timestamp 0
transform 1 0 3220 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _206_
timestamp 0
transform -1 0 4324 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _207_
timestamp 0
transform -1 0 3588 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _208_
timestamp 0
transform -1 0 3220 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _209_
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _210_
timestamp 0
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _211_
timestamp 0
transform -1 0 3588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 0
transform -1 0 6440 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _213_
timestamp 0
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 0
transform -1 0 8096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _215_
timestamp 0
transform -1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _216_
timestamp 0
transform 1 0 9936 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 0
transform -1 0 10304 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _218_
timestamp 0
transform 1 0 10212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _219_
timestamp 0
transform 1 0 10212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _220_
timestamp 0
transform 1 0 7820 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _221_
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _222_
timestamp 0
transform -1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 0
transform -1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _224_
timestamp 0
transform -1 0 4048 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _225_
timestamp 0
transform -1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _226_
timestamp 0
transform 1 0 1748 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _227_
timestamp 0
transform 1 0 2668 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _228_
timestamp 0
transform 1 0 1472 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _229_
timestamp 0
transform 1 0 4324 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _230_
timestamp 0
transform 1 0 4784 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _231_
timestamp 0
transform -1 0 8280 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _232_
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _233_
timestamp 0
transform 1 0 9108 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _235_
timestamp 0
transform 1 0 9016 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _236_
timestamp 0
transform 1 0 9108 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _237_
timestamp 0
transform 1 0 6808 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _238_
timestamp 0
transform 1 0 4968 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _239_
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _240_
timestamp 0
transform 1 0 2024 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 0
transform 1 0 1840 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _242_
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform 1 0 5336 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 0
transform -1 0 4692 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 0
transform 1 0 8004 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_2  clkload0
timestamp 0
transform 1 0 7636 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  clone1
timestamp 0
transform -1 0 4600 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout19
timestamp 0
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout20
timestamp 0
transform 1 0 7176 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout21
timestamp 0
transform -1 0 5888 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout22
timestamp 0
transform -1 0 10764 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23
timestamp 0
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34
timestamp 0
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48
timestamp 0
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52
timestamp 0
transform 1 0 5888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62
timestamp 0
transform 1 0 6808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78
timestamp 0
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 0
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_23
timestamp 0
transform 1 0 3220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_36
timestamp 0
transform 1 0 4416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_43
timestamp 0
transform 1 0 5060 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 0
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_60
timestamp 0
transform 1 0 6624 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_80
timestamp 0
transform 1 0 8464 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_92
timestamp 0
transform 1 0 9568 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_104
timestamp 0
transform 1 0 10672 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_49
timestamp 0
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_59
timestamp 0
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 0
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_105
timestamp 0
transform 1 0 10764 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_11
timestamp 0
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_20
timestamp 0
transform 1 0 2944 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_32
timestamp 0
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 0
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_63
timestamp 0
transform 1 0 6900 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_70
timestamp 0
transform 1 0 7544 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_3_79
timestamp 0
transform 1 0 8372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_88
timestamp 0
transform 1 0 9200 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_96
timestamp 0
transform 1 0 9936 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_100
timestamp 0
transform 1 0 10304 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_58
timestamp 0
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_70
timestamp 0
transform 1 0 7544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_76
timestamp 0
transform 1 0 8096 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 0
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 0
transform 1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_20
timestamp 0
transform 1 0 2944 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_32
timestamp 0
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_41
timestamp 0
transform 1 0 4876 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_45
timestamp 0
transform 1 0 5244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 0
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 0
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 0
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 0
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_36
timestamp 0
transform 1 0 4416 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_60
timestamp 0
transform 1 0 6624 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_90
timestamp 0
transform 1 0 9384 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_105
timestamp 0
transform 1 0 10764 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_7_38
timestamp 0
transform 1 0 4600 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_44
timestamp 0
transform 1 0 5152 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_100
timestamp 0
transform 1 0 10304 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_106
timestamp 0
transform 1 0 10856 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_32
timestamp 0
transform 1 0 4048 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_44
timestamp 0
transform 1 0 5152 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_76
timestamp 0
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 0
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_10
timestamp 0
transform 1 0 2024 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_14
timestamp 0
transform 1 0 2392 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_26
timestamp 0
transform 1 0 3496 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_47
timestamp 0
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 0
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_95
timestamp 0
transform 1 0 9844 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 0
transform 1 0 7452 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_76
timestamp 0
transform 1 0 8096 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_105
timestamp 0
transform 1 0 10764 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 0
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_60
timestamp 0
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_95
timestamp 0
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_102
timestamp 0
transform 1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_106
timestamp 0
transform 1 0 10856 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_23
timestamp 0
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_38
timestamp 0
transform 1 0 4600 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_12_60
timestamp 0
transform 1 0 6624 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 0
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_106
timestamp 0
transform 1 0 10856 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_9
timestamp 0
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_30
timestamp 0
transform 1 0 3864 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_38
timestamp 0
transform 1 0 4600 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 0
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_73
timestamp 0
transform 1 0 7820 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_89
timestamp 0
transform 1 0 9292 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_97
timestamp 0
transform 1 0 10028 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_102
timestamp 0
transform 1 0 10488 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_106
timestamp 0
transform 1 0 10856 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 0
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_37
timestamp 0
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_62
timestamp 0
transform 1 0 6808 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_78
timestamp 0
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_21
timestamp 0
transform 1 0 3036 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 0
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_99
timestamp 0
transform 1 0 10212 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_37
timestamp 0
transform 1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_59
timestamp 0
transform 1 0 6532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_63
timestamp 0
transform 1 0 6900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 0
transform 1 0 7544 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 0
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_98
timestamp 0
transform 1 0 10120 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_106
timestamp 0
transform 1 0 10856 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_29
timestamp 0
transform 1 0 3772 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_34
timestamp 0
transform 1 0 4232 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_42
timestamp 0
transform 1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_48
timestamp 0
transform 1 0 5520 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_65
timestamp 0
transform 1 0 7084 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 0
transform 1 0 8096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_83
timestamp 0
transform 1 0 8740 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_91
timestamp 0
transform 1 0 9476 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_103
timestamp 0
transform 1 0 10580 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform -1 0 3220 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 4508 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 0
transform -1 0 3588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 0
transform -1 0 9476 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 0
transform -1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 0
transform -1 0 5520 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 0
transform -1 0 6164 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 0
transform -1 0 4232 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 0
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 0
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 0
transform 1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 0
transform -1 0 6256 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 0
transform -1 0 8004 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 0
transform -1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 0
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 0
transform -1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 0
transform -1 0 7452 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 0
transform -1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 0
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_18
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 11224 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_19
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_20
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_21
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 11224 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_22
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 11224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_23
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 11224 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_24
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 11224 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_25
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 11224 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_26
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 11224 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_27
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 11224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_28
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_29
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 11224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_30
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_31
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 11224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_32
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_33
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 11224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_34
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 11224 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_35
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 11224 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  rebuffer2
timestamp 0
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer3
timestamp 0
transform -1 0 4508 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_36
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_37
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_39
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_40
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_41
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_42
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_43
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_44
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_45
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_46
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_47
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_48
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_49
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_50
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_51
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_52
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_53
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_54
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_55
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_56
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_57
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_58
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_59
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_60
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_61
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_62
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_63
timestamp 0
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_64
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_65
timestamp 0
transform 1 0 8832 0 -1 11968
box -38 -48 130 592
<< labels >>
rlabel metal1 s 6164 11968 6164 11968 4 VGND
rlabel metal1 s 6164 11424 6164 11424 4 VPWR
rlabel metal1 s 2116 6426 2116 6426 4 _000_
rlabel metal1 s 9614 10098 9614 10098 4 _001_
rlabel metal1 s 7268 7990 7268 7990 4 _002_
rlabel metal2 s 5290 8500 5290 8500 4 _003_
rlabel metal1 s 3726 7310 3726 7310 4 _004_
rlabel metal2 s 2806 9316 2806 9316 4 _005_
rlabel metal2 s 2162 10268 2162 10268 4 _006_
rlabel metal2 s 3082 6052 3082 6052 4 _007_
rlabel metal2 s 1794 4760 1794 4760 4 _008_
rlabel metal1 s 4784 3978 4784 3978 4 _009_
rlabel metal2 s 5106 5916 5106 5916 4 _010_
rlabel metal1 s 7958 6392 7958 6392 4 _011_
rlabel metal1 s 9292 4658 9292 4658 4 _012_
rlabel metal1 s 9246 5134 9246 5134 4 _013_
rlabel metal1 s 9384 6426 9384 6426 4 _014_
rlabel metal2 s 9246 8738 9246 8738 4 _015_
rlabel metal1 s 3595 6698 3595 6698 4 _016_
rlabel metal1 s 3956 5882 3956 5882 4 _017_
rlabel metal1 s 3227 4522 3227 4522 4 _018_
rlabel metal1 s 6079 4522 6079 4522 4 _019_
rlabel metal2 s 5842 6392 5842 6392 4 _020_
rlabel metal2 s 7498 6494 7498 6494 4 _021_
rlabel metal1 s 10074 4114 10074 4114 4 _022_
rlabel metal2 s 10074 5406 10074 5406 4 _023_
rlabel metal1 s 10212 6426 10212 6426 4 _024_
rlabel metal2 s 10350 8738 10350 8738 4 _025_
rlabel metal1 s 10396 9622 10396 9622 4 _026_
rlabel metal1 s 7912 8058 7912 8058 4 _027_
rlabel metal2 s 6394 8058 6394 8058 4 _028_
rlabel metal1 s 4738 8330 4738 8330 4 _029_
rlabel metal1 s 4278 9146 4278 9146 4 _030_
rlabel metal2 s 3910 10200 3910 10200 4 _031_
rlabel metal2 s 3358 7650 3358 7650 4 _032_
rlabel metal1 s 1518 7242 1518 7242 4 _033_
rlabel metal1 s 5382 3468 5382 3468 4 _034_
rlabel metal1 s 4830 3162 4830 3162 4 _035_
rlabel metal1 s 5060 3502 5060 3502 4 _036_
rlabel metal2 s 5566 3876 5566 3876 4 _037_
rlabel metal1 s 7314 4046 7314 4046 4 _038_
rlabel metal1 s 6946 3434 6946 3434 4 _039_
rlabel metal1 s 7222 3094 7222 3094 4 _040_
rlabel metal1 s 7222 2414 7222 2414 4 _041_
rlabel metal1 s 7268 2618 7268 2618 4 _042_
rlabel metal1 s 7544 3706 7544 3706 4 _043_
rlabel metal1 s 7222 2992 7222 2992 4 _044_
rlabel metal1 s 7222 2550 7222 2550 4 _045_
rlabel metal1 s 6716 3706 6716 3706 4 _046_
rlabel metal2 s 7866 3638 7866 3638 4 _047_
rlabel metal1 s 7038 4182 7038 4182 4 _048_
rlabel metal1 s 7084 3910 7084 3910 4 _049_
rlabel metal1 s 7958 10574 7958 10574 4 _050_
rlabel metal1 s 6670 10234 6670 10234 4 _051_
rlabel metal1 s 7636 10574 7636 10574 4 _052_
rlabel metal1 s 6118 8432 6118 8432 4 _053_
rlabel metal1 s 3128 5814 3128 5814 4 _054_
rlabel metal1 s 2898 5576 2898 5576 4 _055_
rlabel metal1 s 2392 4250 2392 4250 4 _056_
rlabel metal1 s 2476 5338 2476 5338 4 _057_
rlabel metal1 s 4784 4250 4784 4250 4 _058_
rlabel metal1 s 7314 5780 7314 5780 4 _059_
rlabel metal1 s 5934 6120 5934 6120 4 _060_
rlabel metal2 s 4646 6120 4646 6120 4 _061_
rlabel metal1 s 7314 5882 7314 5882 4 _062_
rlabel metal1 s 8372 5882 8372 5882 4 _063_
rlabel metal1 s 7728 5882 7728 5882 4 _064_
rlabel metal1 s 8924 5678 8924 5678 4 _065_
rlabel metal1 s 8694 4794 8694 4794 4 _066_
rlabel metal2 s 8878 4760 8878 4760 4 _067_
rlabel metal1 s 8556 5338 8556 5338 4 _068_
rlabel metal1 s 8740 5882 8740 5882 4 _069_
rlabel metal1 s 9660 6358 9660 6358 4 _070_
rlabel metal1 s 8188 8942 8188 8942 4 _071_
rlabel metal1 s 9108 8602 9108 8602 4 _072_
rlabel metal1 s 9016 8330 9016 8330 4 _073_
rlabel metal1 s 9430 9690 9430 9690 4 _074_
rlabel metal1 s 7636 7786 7636 7786 4 _075_
rlabel metal2 s 6578 9146 6578 9146 4 _076_
rlabel metal1 s 5244 8602 5244 8602 4 _077_
rlabel metal1 s 5374 8874 5374 8874 4 _078_
rlabel metal1 s 4324 8942 4324 8942 4 _079_
rlabel metal1 s 3450 7922 3450 7922 4 _080_
rlabel metal1 s 3450 9146 3450 9146 4 _081_
rlabel metal2 s 2982 8874 2982 8874 4 _082_
rlabel metal1 s 4738 10676 4738 10676 4 _083_
rlabel metal2 s 5198 11322 5198 11322 4 _084_
rlabel metal2 s 6210 8262 6210 8262 4 _085_
rlabel metal2 s 5934 10506 5934 10506 4 _086_
rlabel metal1 s 8464 10234 8464 10234 4 _087_
rlabel metal1 s 7544 10982 7544 10982 4 _088_
rlabel metal1 s 8878 4080 8878 4080 4 _089_
rlabel metal1 s 7682 2448 7682 2448 4 _090_
rlabel metal1 s 6302 3162 6302 3162 4 _091_
rlabel metal1 s 5612 3026 5612 3026 4 _092_
rlabel metal1 s 4232 3434 4232 3434 4 _093_
rlabel metal1 s 4094 3060 4094 3060 4 _094_
rlabel metal1 s 3910 3060 3910 3060 4 _095_
rlabel metal2 s 5106 10370 5106 10370 4 _096_
rlabel metal1 s 4922 10098 4922 10098 4 _097_
rlabel metal1 s 5796 10710 5796 10710 4 _098_
rlabel metal2 s 5566 9826 5566 9826 4 _099_
rlabel metal1 s 5566 9486 5566 9486 4 _100_
rlabel metal1 s 6578 10642 6578 10642 4 _101_
rlabel metal1 s 5474 10064 5474 10064 4 _102_
rlabel metal2 s 6578 10234 6578 10234 4 _103_
rlabel metal1 s 9246 11186 9246 11186 4 _104_
rlabel metal2 s 9430 11492 9430 11492 4 _105_
rlabel metal2 s 8418 11526 8418 11526 4 _106_
rlabel metal2 s 7958 10370 7958 10370 4 _107_
rlabel metal2 s 7958 11526 7958 11526 4 _108_
rlabel metal1 s 7314 11118 7314 11118 4 _109_
rlabel metal1 s 8188 10642 8188 10642 4 _110_
rlabel metal1 s 7406 9996 7406 9996 4 _111_
rlabel metal1 s 6854 9962 6854 9962 4 _112_
rlabel metal2 s 5382 8177 5382 8177 4 clk
rlabel metal2 s 6670 7752 6670 7752 4 clknet_0_clk
rlabel metal1 s 1656 6834 1656 6834 4 clknet_1_0__leaf_clk
rlabel metal2 s 9062 9520 9062 9520 4 clknet_1_1__leaf_clk
rlabel metal2 s 3542 2822 3542 2822 4 net1
rlabel metal1 s 5244 2618 5244 2618 4 net10
rlabel metal1 s 6302 2618 6302 2618 4 net11
rlabel metal1 s 8142 2856 8142 2856 4 net12
rlabel metal1 s 7820 2618 7820 2618 4 net13
rlabel metal1 s 8648 2618 8648 2618 4 net14
rlabel metal1 s 8510 11594 8510 11594 4 net15
rlabel metal2 s 7590 10812 7590 10812 4 net16
rlabel metal1 s 10534 5610 10534 5610 4 net17
rlabel metal2 s 3174 8262 3174 8262 4 net18
rlabel metal1 s 2346 6120 2346 6120 4 net19
rlabel metal1 s 9706 11084 9706 11084 4 net2
rlabel metal2 s 10074 9486 10074 9486 4 net20
rlabel metal1 s 4508 8942 4508 8942 4 net21
rlabel metal2 s 10258 9010 10258 9010 4 net22
rlabel metal2 s 2714 9248 2714 9248 4 net23
rlabel metal1 s 3910 9622 3910 9622 4 net24
rlabel metal1 s 3358 8976 3358 8976 4 net25
rlabel metal1 s 2162 7378 2162 7378 4 net26
rlabel metal1 s 3358 10778 3358 10778 4 net27
rlabel metal2 s 8509 11118 8509 11118 4 net3
rlabel metal2 s 6486 11356 6486 11356 4 net4
rlabel metal1 s 6210 11118 6210 11118 4 net5
rlabel metal1 s 4692 11730 4692 11730 4 net6
rlabel metal1 s 4600 10642 4600 10642 4 net7
rlabel metal1 s 4508 2550 4508 2550 4 net8
rlabel metal1 s 4600 3026 4600 3026 4 net9
rlabel metal3 s 1096 7548 1096 7548 4 out
rlabel metal2 s 3266 1588 3266 1588 4 psc[0]
rlabel metal1 s 9154 11730 9154 11730 4 psc[10]
rlabel metal2 s 8418 13105 8418 13105 4 psc[11]
rlabel metal2 s 5244 12716 5244 12716 4 psc[12]
rlabel metal1 s 5888 11730 5888 11730 4 psc[13]
rlabel metal1 s 4738 11798 4738 11798 4 psc[14]
rlabel metal1 s 3956 11730 3956 11730 4 psc[15]
rlabel metal2 s 3910 1588 3910 1588 4 psc[1]
rlabel metal2 s 4554 1588 4554 1588 4 psc[2]
rlabel metal2 s 5198 1027 5198 1027 4 psc[3]
rlabel metal2 s 6486 1520 6486 1520 4 psc[4]
rlabel metal2 s 7130 1520 7130 1520 4 psc[5]
rlabel metal2 s 7774 1588 7774 1588 4 psc[6]
rlabel metal2 s 8418 1588 8418 1588 4 psc[7]
rlabel metal1 s 7820 11730 7820 11730 4 psc[8]
rlabel metal1 s 7176 11730 7176 11730 4 psc[9]
rlabel metal1 s 2346 5712 2346 5712 4 psc_cnt\[0\]
rlabel metal1 s 8142 9656 8142 9656 4 psc_cnt\[10\]
rlabel metal1 s 8924 11118 8924 11118 4 psc_cnt\[11\]
rlabel metal1 s 6394 8908 6394 8908 4 psc_cnt\[12\]
rlabel metal2 s 6026 8194 6026 8194 4 psc_cnt\[13\]
rlabel metal1 s 5336 10642 5336 10642 4 psc_cnt\[14\]
rlabel metal2 s 3542 10438 3542 10438 4 psc_cnt\[15\]
rlabel metal2 s 2714 5440 2714 5440 4 psc_cnt\[1\]
rlabel metal2 s 2530 4964 2530 4964 4 psc_cnt\[2\]
rlabel metal1 s 5474 4114 5474 4114 4 psc_cnt\[3\]
rlabel metal2 s 6563 2414 6563 2414 4 psc_cnt\[4\]
rlabel metal1 s 6945 3026 6945 3026 4 psc_cnt\[5\]
rlabel metal1 s 8418 4488 8418 4488 4 psc_cnt\[6\]
rlabel metal2 s 9154 4556 9154 4556 4 psc_cnt\[7\]
rlabel metal2 s 8326 7106 8326 7106 4 psc_cnt\[8\]
rlabel metal2 s 8234 9860 8234 9860 4 psc_cnt\[9\]
rlabel metal2 s 10902 4471 10902 4471 4 rst
flabel metal4 s 4868 2128 5188 12016 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4208 2128 4528 12016 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 9528 800 9648 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal3 s 0 7488 800 7608 0 FreeSans 600 0 0 0 out
port 4 nsew
flabel metal2 s 3238 0 3294 800 0 FreeSans 280 90 0 0 psc[0]
port 5 nsew
flabel metal2 s 9034 13716 9090 14516 0 FreeSans 280 90 0 0 psc[10]
port 6 nsew
flabel metal2 s 8390 13716 8446 14516 0 FreeSans 280 90 0 0 psc[11]
port 7 nsew
flabel metal2 s 5170 13716 5226 14516 0 FreeSans 280 90 0 0 psc[12]
port 8 nsew
flabel metal2 s 5814 13716 5870 14516 0 FreeSans 280 90 0 0 psc[13]
port 9 nsew
flabel metal2 s 4526 13716 4582 14516 0 FreeSans 280 90 0 0 psc[14]
port 10 nsew
flabel metal2 s 3882 13716 3938 14516 0 FreeSans 280 90 0 0 psc[15]
port 11 nsew
flabel metal2 s 3882 0 3938 800 0 FreeSans 280 90 0 0 psc[1]
port 12 nsew
flabel metal2 s 4526 0 4582 800 0 FreeSans 280 90 0 0 psc[2]
port 13 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 psc[3]
port 14 nsew
flabel metal2 s 6458 0 6514 800 0 FreeSans 280 90 0 0 psc[4]
port 15 nsew
flabel metal2 s 7102 0 7158 800 0 FreeSans 280 90 0 0 psc[5]
port 16 nsew
flabel metal2 s 7746 0 7802 800 0 FreeSans 280 90 0 0 psc[6]
port 17 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 psc[7]
port 18 nsew
flabel metal2 s 7746 13716 7802 14516 0 FreeSans 280 90 0 0 psc[8]
port 19 nsew
flabel metal2 s 7102 13716 7158 14516 0 FreeSans 280 90 0 0 psc[9]
port 20 nsew
flabel metal3 s 11572 4768 12372 4888 0 FreeSans 600 0 0 0 rst
port 21 nsew
<< properties >>
string FIXED_BBOX 0 0 12372 14516
<< end >>
