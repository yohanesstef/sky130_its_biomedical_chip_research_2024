magic
tech sky130A
magscale 1 2
timestamp 1730019635
<< error_p >>
rect 19 207 77 213
rect 19 173 31 207
rect 19 167 77 173
rect -77 -173 -19 -167
rect -77 -207 -65 -173
rect -77 -213 -19 -207
<< nwell >>
rect -65 188 161 226
rect -161 -188 161 188
rect -161 -226 65 -188
<< pmos >>
rect -63 -126 -33 126
rect 33 -126 63 126
<< pdiff >>
rect -125 114 -63 126
rect -125 -114 -113 114
rect -79 -114 -63 114
rect -125 -126 -63 -114
rect -33 114 33 126
rect -33 -114 -17 114
rect 17 -114 33 114
rect -33 -126 33 -114
rect 63 114 125 126
rect 63 -114 79 114
rect 113 -114 125 114
rect 63 -126 125 -114
<< pdiffc >>
rect -113 -114 -79 114
rect -17 -114 17 114
rect 79 -114 113 114
<< poly >>
rect 15 207 81 223
rect 15 173 31 207
rect 65 173 81 207
rect 15 157 81 173
rect -63 126 -33 152
rect 33 126 63 157
rect -63 -157 -33 -126
rect 33 -152 63 -126
rect -81 -173 -15 -157
rect -81 -207 -65 -173
rect -31 -207 -15 -173
rect -81 -223 -15 -207
<< polycont >>
rect 31 173 65 207
rect -65 -207 -31 -173
<< locali >>
rect 15 173 31 207
rect 65 173 81 207
rect -113 114 -79 130
rect -113 -130 -79 -114
rect -17 114 17 130
rect -17 -130 17 -114
rect 79 114 113 130
rect 79 -130 113 -114
rect -81 -207 -65 -173
rect -31 -207 -15 -173
<< viali >>
rect 31 173 65 207
rect -113 -114 -79 114
rect -17 -114 17 114
rect 79 -114 113 114
rect -65 -207 -31 -173
<< metal1 >>
rect 19 207 77 213
rect 19 173 31 207
rect 65 173 77 207
rect 19 167 77 173
rect -119 114 -73 126
rect -119 -114 -113 114
rect -79 -114 -73 114
rect -119 -126 -73 -114
rect -23 114 23 126
rect -23 -114 -17 114
rect 17 -114 23 114
rect -23 -126 23 -114
rect 73 114 119 126
rect 73 -114 79 114
rect 113 -114 119 114
rect 73 -126 119 -114
rect -77 -173 -19 -167
rect -77 -207 -65 -173
rect -31 -207 -19 -173
rect -77 -213 -19 -207
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.26 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
